module  TABLE(exp, value); 
input  [11:0]   exp;   
output [15:0]   value; 
reg    [15:0]   value; 

always @(*)begin   
	 case(exp)   
          'd0000 : value = 'h1000;    //value='d 4096;             
          'd0001 : value = 'h1002;    //value='d 4098;             
          'd0002 : value = 'h1004;    //value='d 4100;             
          'd0003 : value = 'h1006;    //value='d 4102;             
          'd0004 : value = 'h1009;    //value='d 4105;             
          'd0005 : value = 'h100B;    //value='d 4107;             
          'd0006 : value = 'h100D;    //value='d 4109;             
          'd0007 : value = 'h1010;    //value='d 4112;             
          'd0008 : value = 'h1012;    //value='d 4114;             
          'd0009 : value = 'h1014;    //value='d 4116;             
          'd0010 : value = 'h1017;    //value='d 4119;             
          'd0011 : value = 'h1019;    //value='d 4121;             
          'd0012 : value = 'h101B;    //value='d 4123;             
          'd0013 : value = 'h101E;    //value='d 4126;             
          'd0014 : value = 'h1020;    //value='d 4128;             
          'd0015 : value = 'h1022;    //value='d 4130;             
          'd0016 : value = 'h1025;    //value='d 4133;             
          'd0017 : value = 'h1027;    //value='d 4135;             
          'd0018 : value = 'h1029;    //value='d 4137;             
          'd0019 : value = 'h102B;    //value='d 4139;             
          'd0020 : value = 'h102E;    //value='d 4142;             
          'd0021 : value = 'h1030;    //value='d 4144;             
          'd0022 : value = 'h1032;    //value='d 4146;             
          'd0023 : value = 'h1035;    //value='d 4149;             
          'd0024 : value = 'h1037;    //value='d 4151;             
          'd0025 : value = 'h1039;    //value='d 4153;             
          'd0026 : value = 'h103C;    //value='d 4156;             
          'd0027 : value = 'h103E;    //value='d 4158;             
          'd0028 : value = 'h1040;    //value='d 4160;             
          'd0029 : value = 'h1043;    //value='d 4163;             
          'd0030 : value = 'h1045;    //value='d 4165;             
          'd0031 : value = 'h1048;    //value='d 4168;             
          'd0032 : value = 'h104A;    //value='d 4170;             
          'd0033 : value = 'h104C;    //value='d 4172;             
          'd0034 : value = 'h104F;    //value='d 4175;             
          'd0035 : value = 'h1051;    //value='d 4177;             
          'd0036 : value = 'h1053;    //value='d 4179;             
          'd0037 : value = 'h1056;    //value='d 4182;             
          'd0038 : value = 'h1058;    //value='d 4184;             
          'd0039 : value = 'h105A;    //value='d 4186;             
          'd0040 : value = 'h105D;    //value='d 4189;             
          'd0041 : value = 'h105F;    //value='d 4191;             
          'd0042 : value = 'h1061;    //value='d 4193;             
          'd0043 : value = 'h1064;    //value='d 4196;             
          'd0044 : value = 'h1066;    //value='d 4198;             
          'd0045 : value = 'h1068;    //value='d 4200;             
          'd0046 : value = 'h106B;    //value='d 4203;             
          'd0047 : value = 'h106D;    //value='d 4205;             
          'd0048 : value = 'h1070;    //value='d 4208;             
          'd0049 : value = 'h1072;    //value='d 4210;             
          'd0050 : value = 'h1074;    //value='d 4212;             
          'd0051 : value = 'h1077;    //value='d 4215;             
          'd0052 : value = 'h1079;    //value='d 4217;             
          'd0053 : value = 'h107B;    //value='d 4219;             
          'd0054 : value = 'h107E;    //value='d 4222;             
          'd0055 : value = 'h1080;    //value='d 4224;             
          'd0056 : value = 'h1082;    //value='d 4226;             
          'd0057 : value = 'h1085;    //value='d 4229;             
          'd0058 : value = 'h1087;    //value='d 4231;             
          'd0059 : value = 'h108A;    //value='d 4234;             
          'd0060 : value = 'h108C;    //value='d 4236;             
          'd0061 : value = 'h108E;    //value='d 4238;             
          'd0062 : value = 'h1091;    //value='d 4241;             
          'd0063 : value = 'h1093;    //value='d 4243;             
          'd0064 : value = 'h1096;    //value='d 4246;             
          'd0065 : value = 'h1098;    //value='d 4248;             
          'd0066 : value = 'h109A;    //value='d 4250;             
          'd0067 : value = 'h109D;    //value='d 4253;             
          'd0068 : value = 'h109F;    //value='d 4255;             
          'd0069 : value = 'h10A1;    //value='d 4257;             
          'd0070 : value = 'h10A4;    //value='d 4260;             
          'd0071 : value = 'h10A6;    //value='d 4262;             
          'd0072 : value = 'h10A9;    //value='d 4265;             
          'd0073 : value = 'h10AB;    //value='d 4267;             
          'd0074 : value = 'h10AD;    //value='d 4269;             
          'd0075 : value = 'h10B0;    //value='d 4272;             
          'd0076 : value = 'h10B2;    //value='d 4274;             
          'd0077 : value = 'h10B5;    //value='d 4277;             
          'd0078 : value = 'h10B7;    //value='d 4279;             
          'd0079 : value = 'h10BA;    //value='d 4282;             
          'd0080 : value = 'h10BC;    //value='d 4284;             
          'd0081 : value = 'h10BE;    //value='d 4286;             
          'd0082 : value = 'h10C1;    //value='d 4289;             
          'd0083 : value = 'h10C3;    //value='d 4291;             
          'd0084 : value = 'h10C6;    //value='d 4294;             
          'd0085 : value = 'h10C8;    //value='d 4296;             
          'd0086 : value = 'h10CA;    //value='d 4298;             
          'd0087 : value = 'h10CD;    //value='d 4301;             
          'd0088 : value = 'h10CF;    //value='d 4303;             
          'd0089 : value = 'h10D2;    //value='d 4306;             
          'd0090 : value = 'h10D4;    //value='d 4308;             
          'd0091 : value = 'h10D6;    //value='d 4310;             
          'd0092 : value = 'h10D9;    //value='d 4313;             
          'd0093 : value = 'h10DB;    //value='d 4315;             
          'd0094 : value = 'h10DE;    //value='d 4318;             
          'd0095 : value = 'h10E0;    //value='d 4320;             
          'd0096 : value = 'h10E3;    //value='d 4323;             
          'd0097 : value = 'h10E5;    //value='d 4325;             
          'd0098 : value = 'h10E7;    //value='d 4327;             
          'd0099 : value = 'h10EA;    //value='d 4330;             
          'd0100 : value = 'h10EC;    //value='d 4332;             
          'd0101 : value = 'h10EF;    //value='d 4335;             
          'd0102 : value = 'h10F1;    //value='d 4337;             
          'd0103 : value = 'h10F4;    //value='d 4340;             
          'd0104 : value = 'h10F6;    //value='d 4342;             
          'd0105 : value = 'h10F9;    //value='d 4345;             
          'd0106 : value = 'h10FB;    //value='d 4347;             
          'd0107 : value = 'h10FD;    //value='d 4349;             
          'd0108 : value = 'h1100;    //value='d 4352;             
          'd0109 : value = 'h1102;    //value='d 4354;             
          'd0110 : value = 'h1105;    //value='d 4357;             
          'd0111 : value = 'h1107;    //value='d 4359;             
          'd0112 : value = 'h110A;    //value='d 4362;             
          'd0113 : value = 'h110C;    //value='d 4364;             
          'd0114 : value = 'h110F;    //value='d 4367;             
          'd0115 : value = 'h1111;    //value='d 4369;             
          'd0116 : value = 'h1114;    //value='d 4372;             
          'd0117 : value = 'h1116;    //value='d 4374;             
          'd0118 : value = 'h1118;    //value='d 4376;             
          'd0119 : value = 'h111B;    //value='d 4379;             
          'd0120 : value = 'h111D;    //value='d 4381;             
          'd0121 : value = 'h1120;    //value='d 4384;             
          'd0122 : value = 'h1122;    //value='d 4386;             
          'd0123 : value = 'h1125;    //value='d 4389;             
          'd0124 : value = 'h1127;    //value='d 4391;             
          'd0125 : value = 'h112A;    //value='d 4394;             
          'd0126 : value = 'h112C;    //value='d 4396;             
          'd0127 : value = 'h112F;    //value='d 4399;             
          'd0128 : value = 'h1131;    //value='d 4401;             
          'd0129 : value = 'h1134;    //value='d 4404;             
          'd0130 : value = 'h1136;    //value='d 4406;             
          'd0131 : value = 'h1139;    //value='d 4409;             
          'd0132 : value = 'h113B;    //value='d 4411;             
          'd0133 : value = 'h113D;    //value='d 4413;             
          'd0134 : value = 'h1140;    //value='d 4416;             
          'd0135 : value = 'h1142;    //value='d 4418;             
          'd0136 : value = 'h1145;    //value='d 4421;             
          'd0137 : value = 'h1147;    //value='d 4423;             
          'd0138 : value = 'h114A;    //value='d 4426;             
          'd0139 : value = 'h114C;    //value='d 4428;             
          'd0140 : value = 'h114F;    //value='d 4431;             
          'd0141 : value = 'h1151;    //value='d 4433;             
          'd0142 : value = 'h1154;    //value='d 4436;             
          'd0143 : value = 'h1156;    //value='d 4438;             
          'd0144 : value = 'h1159;    //value='d 4441;             
          'd0145 : value = 'h115B;    //value='d 4443;             
          'd0146 : value = 'h115E;    //value='d 4446;             
          'd0147 : value = 'h1160;    //value='d 4448;             
          'd0148 : value = 'h1163;    //value='d 4451;             
          'd0149 : value = 'h1165;    //value='d 4453;             
          'd0150 : value = 'h1168;    //value='d 4456;             
          'd0151 : value = 'h116A;    //value='d 4458;             
          'd0152 : value = 'h116D;    //value='d 4461;             
          'd0153 : value = 'h116F;    //value='d 4463;             
          'd0154 : value = 'h1172;    //value='d 4466;             
          'd0155 : value = 'h1174;    //value='d 4468;             
          'd0156 : value = 'h1177;    //value='d 4471;             
          'd0157 : value = 'h1179;    //value='d 4473;             
          'd0158 : value = 'h117C;    //value='d 4476;             
          'd0159 : value = 'h117E;    //value='d 4478;             
          'd0160 : value = 'h1181;    //value='d 4481;             
          'd0161 : value = 'h1184;    //value='d 4484;             
          'd0162 : value = 'h1186;    //value='d 4486;             
          'd0163 : value = 'h1189;    //value='d 4489;             
          'd0164 : value = 'h118B;    //value='d 4491;             
          'd0165 : value = 'h118E;    //value='d 4494;             
          'd0166 : value = 'h1190;    //value='d 4496;             
          'd0167 : value = 'h1193;    //value='d 4499;             
          'd0168 : value = 'h1195;    //value='d 4501;             
          'd0169 : value = 'h1198;    //value='d 4504;             
          'd0170 : value = 'h119A;    //value='d 4506;             
          'd0171 : value = 'h119D;    //value='d 4509;             
          'd0172 : value = 'h119F;    //value='d 4511;             
          'd0173 : value = 'h11A2;    //value='d 4514;             
          'd0174 : value = 'h11A4;    //value='d 4516;             
          'd0175 : value = 'h11A7;    //value='d 4519;             
          'd0176 : value = 'h11A9;    //value='d 4521;             
          'd0177 : value = 'h11AC;    //value='d 4524;             
          'd0178 : value = 'h11AF;    //value='d 4527;             
          'd0179 : value = 'h11B1;    //value='d 4529;             
          'd0180 : value = 'h11B4;    //value='d 4532;             
          'd0181 : value = 'h11B6;    //value='d 4534;             
          'd0182 : value = 'h11B9;    //value='d 4537;             
          'd0183 : value = 'h11BB;    //value='d 4539;             
          'd0184 : value = 'h11BE;    //value='d 4542;             
          'd0185 : value = 'h11C0;    //value='d 4544;             
          'd0186 : value = 'h11C3;    //value='d 4547;             
          'd0187 : value = 'h11C6;    //value='d 4550;             
          'd0188 : value = 'h11C8;    //value='d 4552;             
          'd0189 : value = 'h11CB;    //value='d 4555;             
          'd0190 : value = 'h11CD;    //value='d 4557;             
          'd0191 : value = 'h11D0;    //value='d 4560;             
          'd0192 : value = 'h11D2;    //value='d 4562;             
          'd0193 : value = 'h11D5;    //value='d 4565;             
          'd0194 : value = 'h11D7;    //value='d 4567;             
          'd0195 : value = 'h11DA;    //value='d 4570;             
          'd0196 : value = 'h11DD;    //value='d 4573;             
          'd0197 : value = 'h11DF;    //value='d 4575;             
          'd0198 : value = 'h11E2;    //value='d 4578;             
          'd0199 : value = 'h11E4;    //value='d 4580;             
          'd0200 : value = 'h11E7;    //value='d 4583;             
          'd0201 : value = 'h11E9;    //value='d 4585;             
          'd0202 : value = 'h11EC;    //value='d 4588;             
          'd0203 : value = 'h11EF;    //value='d 4591;             
          'd0204 : value = 'h11F1;    //value='d 4593;             
          'd0205 : value = 'h11F4;    //value='d 4596;             
          'd0206 : value = 'h11F6;    //value='d 4598;             
          'd0207 : value = 'h11F9;    //value='d 4601;             
          'd0208 : value = 'h11FC;    //value='d 4604;             
          'd0209 : value = 'h11FE;    //value='d 4606;             
          'd0210 : value = 'h1201;    //value='d 4609;             
          'd0211 : value = 'h1203;    //value='d 4611;             
          'd0212 : value = 'h1206;    //value='d 4614;             
          'd0213 : value = 'h1209;    //value='d 4617;             
          'd0214 : value = 'h120B;    //value='d 4619;             
          'd0215 : value = 'h120E;    //value='d 4622;             
          'd0216 : value = 'h1210;    //value='d 4624;             
          'd0217 : value = 'h1213;    //value='d 4627;             
          'd0218 : value = 'h1216;    //value='d 4630;             
          'd0219 : value = 'h1218;    //value='d 4632;             
          'd0220 : value = 'h121B;    //value='d 4635;             
          'd0221 : value = 'h121D;    //value='d 4637;             
          'd0222 : value = 'h1220;    //value='d 4640;             
          'd0223 : value = 'h1223;    //value='d 4643;             
          'd0224 : value = 'h1225;    //value='d 4645;             
          'd0225 : value = 'h1228;    //value='d 4648;             
          'd0226 : value = 'h122A;    //value='d 4650;             
          'd0227 : value = 'h122D;    //value='d 4653;             
          'd0228 : value = 'h1230;    //value='d 4656;             
          'd0229 : value = 'h1232;    //value='d 4658;             
          'd0230 : value = 'h1235;    //value='d 4661;             
          'd0231 : value = 'h1237;    //value='d 4663;             
          'd0232 : value = 'h123A;    //value='d 4666;             
          'd0233 : value = 'h123D;    //value='d 4669;             
          'd0234 : value = 'h123F;    //value='d 4671;             
          'd0235 : value = 'h1242;    //value='d 4674;             
          'd0236 : value = 'h1245;    //value='d 4677;             
          'd0237 : value = 'h1247;    //value='d 4679;             
          'd0238 : value = 'h124A;    //value='d 4682;             
          'd0239 : value = 'h124C;    //value='d 4684;             
          'd0240 : value = 'h124F;    //value='d 4687;             
          'd0241 : value = 'h1252;    //value='d 4690;             
          'd0242 : value = 'h1254;    //value='d 4692;             
          'd0243 : value = 'h1257;    //value='d 4695;             
          'd0244 : value = 'h125A;    //value='d 4698;             
          'd0245 : value = 'h125C;    //value='d 4700;             
          'd0246 : value = 'h125F;    //value='d 4703;             
          'd0247 : value = 'h1262;    //value='d 4706;             
          'd0248 : value = 'h1264;    //value='d 4708;             
          'd0249 : value = 'h1267;    //value='d 4711;             
          'd0250 : value = 'h126A;    //value='d 4714;             
          'd0251 : value = 'h126C;    //value='d 4716;             
          'd0252 : value = 'h126F;    //value='d 4719;             
          'd0253 : value = 'h1272;    //value='d 4722;             
          'd0254 : value = 'h1274;    //value='d 4724;             
          'd0255 : value = 'h1277;    //value='d 4727;             
          'd0256 : value = 'h1279;    //value='d 4729;             
          'd0257 : value = 'h127C;    //value='d 4732;             
          'd0258 : value = 'h127F;    //value='d 4735;             
          'd0259 : value = 'h1281;    //value='d 4737;             
          'd0260 : value = 'h1284;    //value='d 4740;             
          'd0261 : value = 'h1287;    //value='d 4743;             
          'd0262 : value = 'h1289;    //value='d 4745;             
          'd0263 : value = 'h128C;    //value='d 4748;             
          'd0264 : value = 'h128F;    //value='d 4751;             
          'd0265 : value = 'h1291;    //value='d 4753;             
          'd0266 : value = 'h1294;    //value='d 4756;             
          'd0267 : value = 'h1297;    //value='d 4759;             
          'd0268 : value = 'h129A;    //value='d 4762;             
          'd0269 : value = 'h129C;    //value='d 4764;             
          'd0270 : value = 'h129F;    //value='d 4767;             
          'd0271 : value = 'h12A2;    //value='d 4770;             
          'd0272 : value = 'h12A4;    //value='d 4772;             
          'd0273 : value = 'h12A7;    //value='d 4775;             
          'd0274 : value = 'h12AA;    //value='d 4778;             
          'd0275 : value = 'h12AC;    //value='d 4780;             
          'd0276 : value = 'h12AF;    //value='d 4783;             
          'd0277 : value = 'h12B2;    //value='d 4786;             
          'd0278 : value = 'h12B4;    //value='d 4788;             
          'd0279 : value = 'h12B7;    //value='d 4791;             
          'd0280 : value = 'h12BA;    //value='d 4794;             
          'd0281 : value = 'h12BC;    //value='d 4796;             
          'd0282 : value = 'h12BF;    //value='d 4799;             
          'd0283 : value = 'h12C2;    //value='d 4802;             
          'd0284 : value = 'h12C5;    //value='d 4805;             
          'd0285 : value = 'h12C7;    //value='d 4807;             
          'd0286 : value = 'h12CA;    //value='d 4810;             
          'd0287 : value = 'h12CD;    //value='d 4813;             
          'd0288 : value = 'h12CF;    //value='d 4815;             
          'd0289 : value = 'h12D2;    //value='d 4818;             
          'd0290 : value = 'h12D5;    //value='d 4821;             
          'd0291 : value = 'h12D7;    //value='d 4823;             
          'd0292 : value = 'h12DA;    //value='d 4826;             
          'd0293 : value = 'h12DD;    //value='d 4829;             
          'd0294 : value = 'h12E0;    //value='d 4832;             
          'd0295 : value = 'h12E2;    //value='d 4834;             
          'd0296 : value = 'h12E5;    //value='d 4837;             
          'd0297 : value = 'h12E8;    //value='d 4840;             
          'd0298 : value = 'h12EA;    //value='d 4842;             
          'd0299 : value = 'h12ED;    //value='d 4845;             
          'd0300 : value = 'h12F0;    //value='d 4848;             
          'd0301 : value = 'h12F3;    //value='d 4851;             
          'd0302 : value = 'h12F5;    //value='d 4853;             
          'd0303 : value = 'h12F8;    //value='d 4856;             
          'd0304 : value = 'h12FB;    //value='d 4859;             
          'd0305 : value = 'h12FE;    //value='d 4862;             
          'd0306 : value = 'h1300;    //value='d 4864;             
          'd0307 : value = 'h1303;    //value='d 4867;             
          'd0308 : value = 'h1306;    //value='d 4870;             
          'd0309 : value = 'h1309;    //value='d 4873;             
          'd0310 : value = 'h130B;    //value='d 4875;             
          'd0311 : value = 'h130E;    //value='d 4878;             
          'd0312 : value = 'h1311;    //value='d 4881;             
          'd0313 : value = 'h1314;    //value='d 4884;             
          'd0314 : value = 'h1316;    //value='d 4886;             
          'd0315 : value = 'h1319;    //value='d 4889;             
          'd0316 : value = 'h131C;    //value='d 4892;             
          'd0317 : value = 'h131E;    //value='d 4894;             
          'd0318 : value = 'h1321;    //value='d 4897;             
          'd0319 : value = 'h1324;    //value='d 4900;             
          'd0320 : value = 'h1327;    //value='d 4903;             
          'd0321 : value = 'h132A;    //value='d 4906;             
          'd0322 : value = 'h132C;    //value='d 4908;             
          'd0323 : value = 'h132F;    //value='d 4911;             
          'd0324 : value = 'h1332;    //value='d 4914;             
          'd0325 : value = 'h1335;    //value='d 4917;             
          'd0326 : value = 'h1337;    //value='d 4919;             
          'd0327 : value = 'h133A;    //value='d 4922;             
          'd0328 : value = 'h133D;    //value='d 4925;             
          'd0329 : value = 'h1340;    //value='d 4928;             
          'd0330 : value = 'h1342;    //value='d 4930;             
          'd0331 : value = 'h1345;    //value='d 4933;             
          'd0332 : value = 'h1348;    //value='d 4936;             
          'd0333 : value = 'h134B;    //value='d 4939;             
          'd0334 : value = 'h134E;    //value='d 4942;             
          'd0335 : value = 'h1350;    //value='d 4944;             
          'd0336 : value = 'h1353;    //value='d 4947;             
          'd0337 : value = 'h1356;    //value='d 4950;             
          'd0338 : value = 'h1359;    //value='d 4953;             
          'd0339 : value = 'h135B;    //value='d 4955;             
          'd0340 : value = 'h135E;    //value='d 4958;             
          'd0341 : value = 'h1361;    //value='d 4961;             
          'd0342 : value = 'h1364;    //value='d 4964;             
          'd0343 : value = 'h1367;    //value='d 4967;             
          'd0344 : value = 'h1369;    //value='d 4969;             
          'd0345 : value = 'h136C;    //value='d 4972;             
          'd0346 : value = 'h136F;    //value='d 4975;             
          'd0347 : value = 'h1372;    //value='d 4978;             
          'd0348 : value = 'h1375;    //value='d 4981;             
          'd0349 : value = 'h1377;    //value='d 4983;             
          'd0350 : value = 'h137A;    //value='d 4986;             
          'd0351 : value = 'h137D;    //value='d 4989;             
          'd0352 : value = 'h1380;    //value='d 4992;             
          'd0353 : value = 'h1383;    //value='d 4995;             
          'd0354 : value = 'h1385;    //value='d 4997;             
          'd0355 : value = 'h1388;    //value='d 5000;             
          'd0356 : value = 'h138B;    //value='d 5003;             
          'd0357 : value = 'h138E;    //value='d 5006;             
          'd0358 : value = 'h1391;    //value='d 5009;             
          'd0359 : value = 'h1393;    //value='d 5011;             
          'd0360 : value = 'h1396;    //value='d 5014;             
          'd0361 : value = 'h1399;    //value='d 5017;             
          'd0362 : value = 'h139C;    //value='d 5020;             
          'd0363 : value = 'h139F;    //value='d 5023;             
          'd0364 : value = 'h13A2;    //value='d 5026;             
          'd0365 : value = 'h13A4;    //value='d 5028;             
          'd0366 : value = 'h13A7;    //value='d 5031;             
          'd0367 : value = 'h13AA;    //value='d 5034;             
          'd0368 : value = 'h13AD;    //value='d 5037;             
          'd0369 : value = 'h13B0;    //value='d 5040;             
          'd0370 : value = 'h13B3;    //value='d 5043;             
          'd0371 : value = 'h13B5;    //value='d 5045;             
          'd0372 : value = 'h13B8;    //value='d 5048;             
          'd0373 : value = 'h13BB;    //value='d 5051;             
          'd0374 : value = 'h13BE;    //value='d 5054;             
          'd0375 : value = 'h13C1;    //value='d 5057;             
          'd0376 : value = 'h13C4;    //value='d 5060;             
          'd0377 : value = 'h13C6;    //value='d 5062;             
          'd0378 : value = 'h13C9;    //value='d 5065;             
          'd0379 : value = 'h13CC;    //value='d 5068;             
          'd0380 : value = 'h13CF;    //value='d 5071;             
          'd0381 : value = 'h13D2;    //value='d 5074;             
          'd0382 : value = 'h13D5;    //value='d 5077;             
          'd0383 : value = 'h13D8;    //value='d 5080;             
          'd0384 : value = 'h13DA;    //value='d 5082;             
          'd0385 : value = 'h13DD;    //value='d 5085;             
          'd0386 : value = 'h13E0;    //value='d 5088;             
          'd0387 : value = 'h13E3;    //value='d 5091;             
          'd0388 : value = 'h13E6;    //value='d 5094;             
          'd0389 : value = 'h13E9;    //value='d 5097;             
          'd0390 : value = 'h13EC;    //value='d 5100;             
          'd0391 : value = 'h13EE;    //value='d 5102;             
          'd0392 : value = 'h13F1;    //value='d 5105;             
          'd0393 : value = 'h13F4;    //value='d 5108;             
          'd0394 : value = 'h13F7;    //value='d 5111;             
          'd0395 : value = 'h13FA;    //value='d 5114;             
          'd0396 : value = 'h13FD;    //value='d 5117;             
          'd0397 : value = 'h1400;    //value='d 5120;             
          'd0398 : value = 'h1403;    //value='d 5123;             
          'd0399 : value = 'h1405;    //value='d 5125;             
          'd0400 : value = 'h1408;    //value='d 5128;             
          'd0401 : value = 'h140B;    //value='d 5131;             
          'd0402 : value = 'h140E;    //value='d 5134;             
          'd0403 : value = 'h1411;    //value='d 5137;             
          'd0404 : value = 'h1414;    //value='d 5140;             
          'd0405 : value = 'h1417;    //value='d 5143;             
          'd0406 : value = 'h141A;    //value='d 5146;             
          'd0407 : value = 'h141D;    //value='d 5149;             
          'd0408 : value = 'h141F;    //value='d 5151;             
          'd0409 : value = 'h1422;    //value='d 5154;             
          'd0410 : value = 'h1425;    //value='d 5157;             
          'd0411 : value = 'h1428;    //value='d 5160;             
          'd0412 : value = 'h142B;    //value='d 5163;             
          'd0413 : value = 'h142E;    //value='d 5166;             
          'd0414 : value = 'h1431;    //value='d 5169;             
          'd0415 : value = 'h1434;    //value='d 5172;             
          'd0416 : value = 'h1437;    //value='d 5175;             
          'd0417 : value = 'h143A;    //value='d 5178;             
          'd0418 : value = 'h143C;    //value='d 5180;             
          'd0419 : value = 'h143F;    //value='d 5183;             
          'd0420 : value = 'h1442;    //value='d 5186;             
          'd0421 : value = 'h1445;    //value='d 5189;             
          'd0422 : value = 'h1448;    //value='d 5192;             
          'd0423 : value = 'h144B;    //value='d 5195;             
          'd0424 : value = 'h144E;    //value='d 5198;             
          'd0425 : value = 'h1451;    //value='d 5201;             
          'd0426 : value = 'h1454;    //value='d 5204;             
          'd0427 : value = 'h1457;    //value='d 5207;             
          'd0428 : value = 'h145A;    //value='d 5210;             
          'd0429 : value = 'h145D;    //value='d 5213;             
          'd0430 : value = 'h1460;    //value='d 5216;             
          'd0431 : value = 'h1462;    //value='d 5218;             
          'd0432 : value = 'h1465;    //value='d 5221;             
          'd0433 : value = 'h1468;    //value='d 5224;             
          'd0434 : value = 'h146B;    //value='d 5227;             
          'd0435 : value = 'h146E;    //value='d 5230;             
          'd0436 : value = 'h1471;    //value='d 5233;             
          'd0437 : value = 'h1474;    //value='d 5236;             
          'd0438 : value = 'h1477;    //value='d 5239;             
          'd0439 : value = 'h147A;    //value='d 5242;             
          'd0440 : value = 'h147D;    //value='d 5245;             
          'd0441 : value = 'h1480;    //value='d 5248;             
          'd0442 : value = 'h1483;    //value='d 5251;             
          'd0443 : value = 'h1486;    //value='d 5254;             
          'd0444 : value = 'h1489;    //value='d 5257;             
          'd0445 : value = 'h148C;    //value='d 5260;             
          'd0446 : value = 'h148F;    //value='d 5263;             
          'd0447 : value = 'h1492;    //value='d 5266;             
          'd0448 : value = 'h1495;    //value='d 5269;             
          'd0449 : value = 'h1498;    //value='d 5272;             
          'd0450 : value = 'h149B;    //value='d 5275;             
          'd0451 : value = 'h149D;    //value='d 5277;             
          'd0452 : value = 'h14A0;    //value='d 5280;             
          'd0453 : value = 'h14A3;    //value='d 5283;             
          'd0454 : value = 'h14A6;    //value='d 5286;             
          'd0455 : value = 'h14A9;    //value='d 5289;             
          'd0456 : value = 'h14AC;    //value='d 5292;             
          'd0457 : value = 'h14AF;    //value='d 5295;             
          'd0458 : value = 'h14B2;    //value='d 5298;             
          'd0459 : value = 'h14B5;    //value='d 5301;             
          'd0460 : value = 'h14B8;    //value='d 5304;             
          'd0461 : value = 'h14BB;    //value='d 5307;             
          'd0462 : value = 'h14BE;    //value='d 5310;             
          'd0463 : value = 'h14C1;    //value='d 5313;             
          'd0464 : value = 'h14C4;    //value='d 5316;             
          'd0465 : value = 'h14C7;    //value='d 5319;             
          'd0466 : value = 'h14CA;    //value='d 5322;             
          'd0467 : value = 'h14CD;    //value='d 5325;             
          'd0468 : value = 'h14D0;    //value='d 5328;             
          'd0469 : value = 'h14D3;    //value='d 5331;             
          'd0470 : value = 'h14D6;    //value='d 5334;             
          'd0471 : value = 'h14D9;    //value='d 5337;             
          'd0472 : value = 'h14DC;    //value='d 5340;             
          'd0473 : value = 'h14DF;    //value='d 5343;             
          'd0474 : value = 'h14E2;    //value='d 5346;             
          'd0475 : value = 'h14E5;    //value='d 5349;             
          'd0476 : value = 'h14E8;    //value='d 5352;             
          'd0477 : value = 'h14EB;    //value='d 5355;             
          'd0478 : value = 'h14EE;    //value='d 5358;             
          'd0479 : value = 'h14F1;    //value='d 5361;             
          'd0480 : value = 'h14F4;    //value='d 5364;             
          'd0481 : value = 'h14F7;    //value='d 5367;             
          'd0482 : value = 'h14FA;    //value='d 5370;             
          'd0483 : value = 'h14FD;    //value='d 5373;             
          'd0484 : value = 'h1500;    //value='d 5376;             
          'd0485 : value = 'h1503;    //value='d 5379;             
          'd0486 : value = 'h1506;    //value='d 5382;             
          'd0487 : value = 'h1509;    //value='d 5385;             
          'd0488 : value = 'h150C;    //value='d 5388;             
          'd0489 : value = 'h150F;    //value='d 5391;             
          'd0490 : value = 'h1512;    //value='d 5394;             
          'd0491 : value = 'h1516;    //value='d 5398;             
          'd0492 : value = 'h1519;    //value='d 5401;             
          'd0493 : value = 'h151C;    //value='d 5404;             
          'd0494 : value = 'h151F;    //value='d 5407;             
          'd0495 : value = 'h1522;    //value='d 5410;             
          'd0496 : value = 'h1525;    //value='d 5413;             
          'd0497 : value = 'h1528;    //value='d 5416;             
          'd0498 : value = 'h152B;    //value='d 5419;             
          'd0499 : value = 'h152E;    //value='d 5422;             
          'd0500 : value = 'h1531;    //value='d 5425;             
          'd0501 : value = 'h1534;    //value='d 5428;             
          'd0502 : value = 'h1537;    //value='d 5431;             
          'd0503 : value = 'h153A;    //value='d 5434;             
          'd0504 : value = 'h153D;    //value='d 5437;             
          'd0505 : value = 'h1540;    //value='d 5440;             
          'd0506 : value = 'h1543;    //value='d 5443;             
          'd0507 : value = 'h1546;    //value='d 5446;             
          'd0508 : value = 'h1549;    //value='d 5449;             
          'd0509 : value = 'h154C;    //value='d 5452;             
          'd0510 : value = 'h154F;    //value='d 5455;             
          'd0511 : value = 'h1553;    //value='d 5459;             
          'd0512 : value = 'h1556;    //value='d 5462;             
          'd0513 : value = 'h1559;    //value='d 5465;             
          'd0514 : value = 'h155C;    //value='d 5468;             
          'd0515 : value = 'h155F;    //value='d 5471;             
          'd0516 : value = 'h1562;    //value='d 5474;             
          'd0517 : value = 'h1565;    //value='d 5477;             
          'd0518 : value = 'h1568;    //value='d 5480;             
          'd0519 : value = 'h156B;    //value='d 5483;             
          'd0520 : value = 'h156E;    //value='d 5486;             
          'd0521 : value = 'h1571;    //value='d 5489;             
          'd0522 : value = 'h1574;    //value='d 5492;             
          'd0523 : value = 'h1577;    //value='d 5495;             
          'd0524 : value = 'h157B;    //value='d 5499;             
          'd0525 : value = 'h157E;    //value='d 5502;             
          'd0526 : value = 'h1581;    //value='d 5505;             
          'd0527 : value = 'h1584;    //value='d 5508;             
          'd0528 : value = 'h1587;    //value='d 5511;             
          'd0529 : value = 'h158A;    //value='d 5514;             
          'd0530 : value = 'h158D;    //value='d 5517;             
          'd0531 : value = 'h1590;    //value='d 5520;             
          'd0532 : value = 'h1593;    //value='d 5523;             
          'd0533 : value = 'h1596;    //value='d 5526;             
          'd0534 : value = 'h159A;    //value='d 5530;             
          'd0535 : value = 'h159D;    //value='d 5533;             
          'd0536 : value = 'h15A0;    //value='d 5536;             
          'd0537 : value = 'h15A3;    //value='d 5539;             
          'd0538 : value = 'h15A6;    //value='d 5542;             
          'd0539 : value = 'h15A9;    //value='d 5545;             
          'd0540 : value = 'h15AC;    //value='d 5548;             
          'd0541 : value = 'h15AF;    //value='d 5551;             
          'd0542 : value = 'h15B3;    //value='d 5555;             
          'd0543 : value = 'h15B6;    //value='d 5558;             
          'd0544 : value = 'h15B9;    //value='d 5561;             
          'd0545 : value = 'h15BC;    //value='d 5564;             
          'd0546 : value = 'h15BF;    //value='d 5567;             
          'd0547 : value = 'h15C2;    //value='d 5570;             
          'd0548 : value = 'h15C5;    //value='d 5573;             
          'd0549 : value = 'h15C8;    //value='d 5576;             
          'd0550 : value = 'h15CC;    //value='d 5580;             
          'd0551 : value = 'h15CF;    //value='d 5583;             
          'd0552 : value = 'h15D2;    //value='d 5586;             
          'd0553 : value = 'h15D5;    //value='d 5589;             
          'd0554 : value = 'h15D8;    //value='d 5592;             
          'd0555 : value = 'h15DB;    //value='d 5595;             
          'd0556 : value = 'h15DE;    //value='d 5598;             
          'd0557 : value = 'h15E2;    //value='d 5602;             
          'd0558 : value = 'h15E5;    //value='d 5605;             
          'd0559 : value = 'h15E8;    //value='d 5608;             
          'd0560 : value = 'h15EB;    //value='d 5611;             
          'd0561 : value = 'h15EE;    //value='d 5614;             
          'd0562 : value = 'h15F1;    //value='d 5617;             
          'd0563 : value = 'h15F4;    //value='d 5620;             
          'd0564 : value = 'h15F8;    //value='d 5624;             
          'd0565 : value = 'h15FB;    //value='d 5627;             
          'd0566 : value = 'h15FE;    //value='d 5630;             
          'd0567 : value = 'h1601;    //value='d 5633;             
          'd0568 : value = 'h1604;    //value='d 5636;             
          'd0569 : value = 'h1607;    //value='d 5639;             
          'd0570 : value = 'h160B;    //value='d 5643;             
          'd0571 : value = 'h160E;    //value='d 5646;             
          'd0572 : value = 'h1611;    //value='d 5649;             
          'd0573 : value = 'h1614;    //value='d 5652;             
          'd0574 : value = 'h1617;    //value='d 5655;             
          'd0575 : value = 'h161B;    //value='d 5659;             
          'd0576 : value = 'h161E;    //value='d 5662;             
          'd0577 : value = 'h1621;    //value='d 5665;             
          'd0578 : value = 'h1624;    //value='d 5668;             
          'd0579 : value = 'h1627;    //value='d 5671;             
          'd0580 : value = 'h162A;    //value='d 5674;             
          'd0581 : value = 'h162E;    //value='d 5678;             
          'd0582 : value = 'h1631;    //value='d 5681;             
          'd0583 : value = 'h1634;    //value='d 5684;             
          'd0584 : value = 'h1637;    //value='d 5687;             
          'd0585 : value = 'h163A;    //value='d 5690;             
          'd0586 : value = 'h163E;    //value='d 5694;             
          'd0587 : value = 'h1641;    //value='d 5697;             
          'd0588 : value = 'h1644;    //value='d 5700;             
          'd0589 : value = 'h1647;    //value='d 5703;             
          'd0590 : value = 'h164A;    //value='d 5706;             
          'd0591 : value = 'h164E;    //value='d 5710;             
          'd0592 : value = 'h1651;    //value='d 5713;             
          'd0593 : value = 'h1654;    //value='d 5716;             
          'd0594 : value = 'h1657;    //value='d 5719;             
          'd0595 : value = 'h165A;    //value='d 5722;             
          'd0596 : value = 'h165E;    //value='d 5726;             
          'd0597 : value = 'h1661;    //value='d 5729;             
          'd0598 : value = 'h1664;    //value='d 5732;             
          'd0599 : value = 'h1667;    //value='d 5735;             
          'd0600 : value = 'h166B;    //value='d 5739;             
          'd0601 : value = 'h166E;    //value='d 5742;             
          'd0602 : value = 'h1671;    //value='d 5745;             
          'd0603 : value = 'h1674;    //value='d 5748;             
          'd0604 : value = 'h1678;    //value='d 5752;             
          'd0605 : value = 'h167B;    //value='d 5755;             
          'd0606 : value = 'h167E;    //value='d 5758;             
          'd0607 : value = 'h1681;    //value='d 5761;             
          'd0608 : value = 'h1684;    //value='d 5764;             
          'd0609 : value = 'h1688;    //value='d 5768;             
          'd0610 : value = 'h168B;    //value='d 5771;             
          'd0611 : value = 'h168E;    //value='d 5774;             
          'd0612 : value = 'h1691;    //value='d 5777;             
          'd0613 : value = 'h1695;    //value='d 5781;             
          'd0614 : value = 'h1698;    //value='d 5784;             
          'd0615 : value = 'h169B;    //value='d 5787;             
          'd0616 : value = 'h169E;    //value='d 5790;             
          'd0617 : value = 'h16A2;    //value='d 5794;             
          'd0618 : value = 'h16A5;    //value='d 5797;             
          'd0619 : value = 'h16A8;    //value='d 5800;             
          'd0620 : value = 'h16AB;    //value='d 5803;             
          'd0621 : value = 'h16AF;    //value='d 5807;             
          'd0622 : value = 'h16B2;    //value='d 5810;             
          'd0623 : value = 'h16B5;    //value='d 5813;             
          'd0624 : value = 'h16B9;    //value='d 5817;             
          'd0625 : value = 'h16BC;    //value='d 5820;             
          'd0626 : value = 'h16BF;    //value='d 5823;             
          'd0627 : value = 'h16C2;    //value='d 5826;             
          'd0628 : value = 'h16C6;    //value='d 5830;             
          'd0629 : value = 'h16C9;    //value='d 5833;             
          'd0630 : value = 'h16CC;    //value='d 5836;             
          'd0631 : value = 'h16CF;    //value='d 5839;             
          'd0632 : value = 'h16D3;    //value='d 5843;             
          'd0633 : value = 'h16D6;    //value='d 5846;             
          'd0634 : value = 'h16D9;    //value='d 5849;             
          'd0635 : value = 'h16DD;    //value='d 5853;             
          'd0636 : value = 'h16E0;    //value='d 5856;             
          'd0637 : value = 'h16E3;    //value='d 5859;             
          'd0638 : value = 'h16E7;    //value='d 5863;             
          'd0639 : value = 'h16EA;    //value='d 5866;             
          'd0640 : value = 'h16ED;    //value='d 5869;             
          'd0641 : value = 'h16F0;    //value='d 5872;             
          'd0642 : value = 'h16F4;    //value='d 5876;             
          'd0643 : value = 'h16F7;    //value='d 5879;             
          'd0644 : value = 'h16FA;    //value='d 5882;             
          'd0645 : value = 'h16FE;    //value='d 5886;             
          'd0646 : value = 'h1701;    //value='d 5889;             
          'd0647 : value = 'h1704;    //value='d 5892;             
          'd0648 : value = 'h1708;    //value='d 5896;             
          'd0649 : value = 'h170B;    //value='d 5899;             
          'd0650 : value = 'h170E;    //value='d 5902;             
          'd0651 : value = 'h1712;    //value='d 5906;             
          'd0652 : value = 'h1715;    //value='d 5909;             
          'd0653 : value = 'h1718;    //value='d 5912;             
          'd0654 : value = 'h171B;    //value='d 5915;             
          'd0655 : value = 'h171F;    //value='d 5919;             
          'd0656 : value = 'h1722;    //value='d 5922;             
          'd0657 : value = 'h1725;    //value='d 5925;             
          'd0658 : value = 'h1729;    //value='d 5929;             
          'd0659 : value = 'h172C;    //value='d 5932;             
          'd0660 : value = 'h172F;    //value='d 5935;             
          'd0661 : value = 'h1733;    //value='d 5939;             
          'd0662 : value = 'h1736;    //value='d 5942;             
          'd0663 : value = 'h173A;    //value='d 5946;             
          'd0664 : value = 'h173D;    //value='d 5949;             
          'd0665 : value = 'h1740;    //value='d 5952;             
          'd0666 : value = 'h1744;    //value='d 5956;             
          'd0667 : value = 'h1747;    //value='d 5959;             
          'd0668 : value = 'h174A;    //value='d 5962;             
          'd0669 : value = 'h174E;    //value='d 5966;             
          'd0670 : value = 'h1751;    //value='d 5969;             
          'd0671 : value = 'h1754;    //value='d 5972;             
          'd0672 : value = 'h1758;    //value='d 5976;             
          'd0673 : value = 'h175B;    //value='d 5979;             
          'd0674 : value = 'h175E;    //value='d 5982;             
          'd0675 : value = 'h1762;    //value='d 5986;             
          'd0676 : value = 'h1765;    //value='d 5989;             
          'd0677 : value = 'h1768;    //value='d 5992;             
          'd0678 : value = 'h176C;    //value='d 5996;             
          'd0679 : value = 'h176F;    //value='d 5999;             
          'd0680 : value = 'h1773;    //value='d 6003;             
          'd0681 : value = 'h1776;    //value='d 6006;             
          'd0682 : value = 'h1779;    //value='d 6009;             
          'd0683 : value = 'h177D;    //value='d 6013;             
          'd0684 : value = 'h1780;    //value='d 6016;             
          'd0685 : value = 'h1783;    //value='d 6019;             
          'd0686 : value = 'h1787;    //value='d 6023;             
          'd0687 : value = 'h178A;    //value='d 6026;             
          'd0688 : value = 'h178E;    //value='d 6030;             
          'd0689 : value = 'h1791;    //value='d 6033;             
          'd0690 : value = 'h1794;    //value='d 6036;             
          'd0691 : value = 'h1798;    //value='d 6040;             
          'd0692 : value = 'h179B;    //value='d 6043;             
          'd0693 : value = 'h179F;    //value='d 6047;             
          'd0694 : value = 'h17A2;    //value='d 6050;             
          'd0695 : value = 'h17A5;    //value='d 6053;             
          'd0696 : value = 'h17A9;    //value='d 6057;             
          'd0697 : value = 'h17AC;    //value='d 6060;             
          'd0698 : value = 'h17B0;    //value='d 6064;             
          'd0699 : value = 'h17B3;    //value='d 6067;             
          'd0700 : value = 'h17B6;    //value='d 6070;             
          'd0701 : value = 'h17BA;    //value='d 6074;             
          'd0702 : value = 'h17BD;    //value='d 6077;             
          'd0703 : value = 'h17C1;    //value='d 6081;             
          'd0704 : value = 'h17C4;    //value='d 6084;             
          'd0705 : value = 'h17C8;    //value='d 6088;             
          'd0706 : value = 'h17CB;    //value='d 6091;             
          'd0707 : value = 'h17CE;    //value='d 6094;             
          'd0708 : value = 'h17D2;    //value='d 6098;             
          'd0709 : value = 'h17D5;    //value='d 6101;             
          'd0710 : value = 'h17D9;    //value='d 6105;             
          'd0711 : value = 'h17DC;    //value='d 6108;             
          'd0712 : value = 'h17E0;    //value='d 6112;             
          'd0713 : value = 'h17E3;    //value='d 6115;             
          'd0714 : value = 'h17E6;    //value='d 6118;             
          'd0715 : value = 'h17EA;    //value='d 6122;             
          'd0716 : value = 'h17ED;    //value='d 6125;             
          'd0717 : value = 'h17F1;    //value='d 6129;             
          'd0718 : value = 'h17F4;    //value='d 6132;             
          'd0719 : value = 'h17F8;    //value='d 6136;             
          'd0720 : value = 'h17FB;    //value='d 6139;             
          'd0721 : value = 'h17FF;    //value='d 6143;             
          'd0722 : value = 'h1802;    //value='d 6146;             
          'd0723 : value = 'h1805;    //value='d 6149;             
          'd0724 : value = 'h1809;    //value='d 6153;             
          'd0725 : value = 'h180C;    //value='d 6156;             
          'd0726 : value = 'h1810;    //value='d 6160;             
          'd0727 : value = 'h1813;    //value='d 6163;             
          'd0728 : value = 'h1817;    //value='d 6167;             
          'd0729 : value = 'h181A;    //value='d 6170;             
          'd0730 : value = 'h181E;    //value='d 6174;             
          'd0731 : value = 'h1821;    //value='d 6177;             
          'd0732 : value = 'h1825;    //value='d 6181;             
          'd0733 : value = 'h1828;    //value='d 6184;             
          'd0734 : value = 'h182C;    //value='d 6188;             
          'd0735 : value = 'h182F;    //value='d 6191;             
          'd0736 : value = 'h1833;    //value='d 6195;             
          'd0737 : value = 'h1836;    //value='d 6198;             
          'd0738 : value = 'h183A;    //value='d 6202;             
          'd0739 : value = 'h183D;    //value='d 6205;             
          'd0740 : value = 'h1841;    //value='d 6209;             
          'd0741 : value = 'h1844;    //value='d 6212;             
          'd0742 : value = 'h1848;    //value='d 6216;             
          'd0743 : value = 'h184B;    //value='d 6219;             
          'd0744 : value = 'h184F;    //value='d 6223;             
          'd0745 : value = 'h1852;    //value='d 6226;             
          'd0746 : value = 'h1856;    //value='d 6230;             
          'd0747 : value = 'h1859;    //value='d 6233;             
          'd0748 : value = 'h185D;    //value='d 6237;             
          'd0749 : value = 'h1860;    //value='d 6240;             
          'd0750 : value = 'h1864;    //value='d 6244;             
          'd0751 : value = 'h1867;    //value='d 6247;             
          'd0752 : value = 'h186B;    //value='d 6251;             
          'd0753 : value = 'h186E;    //value='d 6254;             
          'd0754 : value = 'h1872;    //value='d 6258;             
          'd0755 : value = 'h1875;    //value='d 6261;             
          'd0756 : value = 'h1879;    //value='d 6265;             
          'd0757 : value = 'h187C;    //value='d 6268;             
          'd0758 : value = 'h1880;    //value='d 6272;             
          'd0759 : value = 'h1883;    //value='d 6275;             
          'd0760 : value = 'h1887;    //value='d 6279;             
          'd0761 : value = 'h188A;    //value='d 6282;             
          'd0762 : value = 'h188E;    //value='d 6286;             
          'd0763 : value = 'h1891;    //value='d 6289;             
          'd0764 : value = 'h1895;    //value='d 6293;             
          'd0765 : value = 'h1898;    //value='d 6296;             
          'd0766 : value = 'h189C;    //value='d 6300;             
          'd0767 : value = 'h189F;    //value='d 6303;             
          'd0768 : value = 'h18A3;    //value='d 6307;             
          'd0769 : value = 'h18A7;    //value='d 6311;             
          'd0770 : value = 'h18AA;    //value='d 6314;             
          'd0771 : value = 'h18AE;    //value='d 6318;             
          'd0772 : value = 'h18B1;    //value='d 6321;             
          'd0773 : value = 'h18B5;    //value='d 6325;             
          'd0774 : value = 'h18B8;    //value='d 6328;             
          'd0775 : value = 'h18BC;    //value='d 6332;             
          'd0776 : value = 'h18BF;    //value='d 6335;             
          'd0777 : value = 'h18C3;    //value='d 6339;             
          'd0778 : value = 'h18C7;    //value='d 6343;             
          'd0779 : value = 'h18CA;    //value='d 6346;             
          'd0780 : value = 'h18CE;    //value='d 6350;             
          'd0781 : value = 'h18D1;    //value='d 6353;             
          'd0782 : value = 'h18D5;    //value='d 6357;             
          'd0783 : value = 'h18D8;    //value='d 6360;             
          'd0784 : value = 'h18DC;    //value='d 6364;             
          'd0785 : value = 'h18E0;    //value='d 6368;             
          'd0786 : value = 'h18E3;    //value='d 6371;             
          'd0787 : value = 'h18E7;    //value='d 6375;             
          'd0788 : value = 'h18EA;    //value='d 6378;             
          'd0789 : value = 'h18EE;    //value='d 6382;             
          'd0790 : value = 'h18F2;    //value='d 6386;             
          'd0791 : value = 'h18F5;    //value='d 6389;             
          'd0792 : value = 'h18F9;    //value='d 6393;             
          'd0793 : value = 'h18FC;    //value='d 6396;             
          'd0794 : value = 'h1900;    //value='d 6400;             
          'd0795 : value = 'h1904;    //value='d 6404;             
          'd0796 : value = 'h1907;    //value='d 6407;             
          'd0797 : value = 'h190B;    //value='d 6411;             
          'd0798 : value = 'h190E;    //value='d 6414;             
          'd0799 : value = 'h1912;    //value='d 6418;             
          'd0800 : value = 'h1916;    //value='d 6422;             
          'd0801 : value = 'h1919;    //value='d 6425;             
          'd0802 : value = 'h191D;    //value='d 6429;             
          'd0803 : value = 'h1920;    //value='d 6432;             
          'd0804 : value = 'h1924;    //value='d 6436;             
          'd0805 : value = 'h1928;    //value='d 6440;             
          'd0806 : value = 'h192B;    //value='d 6443;             
          'd0807 : value = 'h192F;    //value='d 6447;             
          'd0808 : value = 'h1932;    //value='d 6450;             
          'd0809 : value = 'h1936;    //value='d 6454;             
          'd0810 : value = 'h193A;    //value='d 6458;             
          'd0811 : value = 'h193D;    //value='d 6461;             
          'd0812 : value = 'h1941;    //value='d 6465;             
          'd0813 : value = 'h1945;    //value='d 6469;             
          'd0814 : value = 'h1948;    //value='d 6472;             
          'd0815 : value = 'h194C;    //value='d 6476;             
          'd0816 : value = 'h1950;    //value='d 6480;             
          'd0817 : value = 'h1953;    //value='d 6483;             
          'd0818 : value = 'h1957;    //value='d 6487;             
          'd0819 : value = 'h195A;    //value='d 6490;             
          'd0820 : value = 'h195E;    //value='d 6494;             
          'd0821 : value = 'h1962;    //value='d 6498;             
          'd0822 : value = 'h1965;    //value='d 6501;             
          'd0823 : value = 'h1969;    //value='d 6505;             
          'd0824 : value = 'h196D;    //value='d 6509;             
          'd0825 : value = 'h1970;    //value='d 6512;             
          'd0826 : value = 'h1974;    //value='d 6516;             
          'd0827 : value = 'h1978;    //value='d 6520;             
          'd0828 : value = 'h197B;    //value='d 6523;             
          'd0829 : value = 'h197F;    //value='d 6527;             
          'd0830 : value = 'h1983;    //value='d 6531;             
          'd0831 : value = 'h1986;    //value='d 6534;             
          'd0832 : value = 'h198A;    //value='d 6538;             
          'd0833 : value = 'h198E;    //value='d 6542;             
          'd0834 : value = 'h1991;    //value='d 6545;             
          'd0835 : value = 'h1995;    //value='d 6549;             
          'd0836 : value = 'h1999;    //value='d 6553;             
          'd0837 : value = 'h199D;    //value='d 6557;             
          'd0838 : value = 'h19A0;    //value='d 6560;             
          'd0839 : value = 'h19A4;    //value='d 6564;             
          'd0840 : value = 'h19A8;    //value='d 6568;             
          'd0841 : value = 'h19AB;    //value='d 6571;             
          'd0842 : value = 'h19AF;    //value='d 6575;             
          'd0843 : value = 'h19B3;    //value='d 6579;             
          'd0844 : value = 'h19B6;    //value='d 6582;             
          'd0845 : value = 'h19BA;    //value='d 6586;             
          'd0846 : value = 'h19BE;    //value='d 6590;             
          'd0847 : value = 'h19C1;    //value='d 6593;             
          'd0848 : value = 'h19C5;    //value='d 6597;             
          'd0849 : value = 'h19C9;    //value='d 6601;             
          'd0850 : value = 'h19CD;    //value='d 6605;             
          'd0851 : value = 'h19D0;    //value='d 6608;             
          'd0852 : value = 'h19D4;    //value='d 6612;             
          'd0853 : value = 'h19D8;    //value='d 6616;             
          'd0854 : value = 'h19DB;    //value='d 6619;             
          'd0855 : value = 'h19DF;    //value='d 6623;             
          'd0856 : value = 'h19E3;    //value='d 6627;             
          'd0857 : value = 'h19E7;    //value='d 6631;             
          'd0858 : value = 'h19EA;    //value='d 6634;             
          'd0859 : value = 'h19EE;    //value='d 6638;             
          'd0860 : value = 'h19F2;    //value='d 6642;             
          'd0861 : value = 'h19F6;    //value='d 6646;             
          'd0862 : value = 'h19F9;    //value='d 6649;             
          'd0863 : value = 'h19FD;    //value='d 6653;             
          'd0864 : value = 'h1A01;    //value='d 6657;             
          'd0865 : value = 'h1A05;    //value='d 6661;             
          'd0866 : value = 'h1A08;    //value='d 6664;             
          'd0867 : value = 'h1A0C;    //value='d 6668;             
          'd0868 : value = 'h1A10;    //value='d 6672;             
          'd0869 : value = 'h1A14;    //value='d 6676;             
          'd0870 : value = 'h1A17;    //value='d 6679;             
          'd0871 : value = 'h1A1B;    //value='d 6683;             
          'd0872 : value = 'h1A1F;    //value='d 6687;             
          'd0873 : value = 'h1A23;    //value='d 6691;             
          'd0874 : value = 'h1A26;    //value='d 6694;             
          'd0875 : value = 'h1A2A;    //value='d 6698;             
          'd0876 : value = 'h1A2E;    //value='d 6702;             
          'd0877 : value = 'h1A32;    //value='d 6706;             
          'd0878 : value = 'h1A35;    //value='d 6709;             
          'd0879 : value = 'h1A39;    //value='d 6713;             
          'd0880 : value = 'h1A3D;    //value='d 6717;             
          'd0881 : value = 'h1A41;    //value='d 6721;             
          'd0882 : value = 'h1A44;    //value='d 6724;             
          'd0883 : value = 'h1A48;    //value='d 6728;             
          'd0884 : value = 'h1A4C;    //value='d 6732;             
          'd0885 : value = 'h1A50;    //value='d 6736;             
          'd0886 : value = 'h1A54;    //value='d 6740;             
          'd0887 : value = 'h1A57;    //value='d 6743;             
          'd0888 : value = 'h1A5B;    //value='d 6747;             
          'd0889 : value = 'h1A5F;    //value='d 6751;             
          'd0890 : value = 'h1A63;    //value='d 6755;             
          'd0891 : value = 'h1A67;    //value='d 6759;             
          'd0892 : value = 'h1A6A;    //value='d 6762;             
          'd0893 : value = 'h1A6E;    //value='d 6766;             
          'd0894 : value = 'h1A72;    //value='d 6770;             
          'd0895 : value = 'h1A76;    //value='d 6774;             
          'd0896 : value = 'h1A7A;    //value='d 6778;             
          'd0897 : value = 'h1A7D;    //value='d 6781;             
          'd0898 : value = 'h1A81;    //value='d 6785;             
          'd0899 : value = 'h1A85;    //value='d 6789;             
          'd0900 : value = 'h1A89;    //value='d 6793;             
          'd0901 : value = 'h1A8D;    //value='d 6797;             
          'd0902 : value = 'h1A91;    //value='d 6801;             
          'd0903 : value = 'h1A94;    //value='d 6804;             
          'd0904 : value = 'h1A98;    //value='d 6808;             
          'd0905 : value = 'h1A9C;    //value='d 6812;             
          'd0906 : value = 'h1AA0;    //value='d 6816;             
          'd0907 : value = 'h1AA4;    //value='d 6820;             
          'd0908 : value = 'h1AA8;    //value='d 6824;             
          'd0909 : value = 'h1AAB;    //value='d 6827;             
          'd0910 : value = 'h1AAF;    //value='d 6831;             
          'd0911 : value = 'h1AB3;    //value='d 6835;             
          'd0912 : value = 'h1AB7;    //value='d 6839;             
          'd0913 : value = 'h1ABB;    //value='d 6843;             
          'd0914 : value = 'h1ABF;    //value='d 6847;             
          'd0915 : value = 'h1AC2;    //value='d 6850;             
          'd0916 : value = 'h1AC6;    //value='d 6854;             
          'd0917 : value = 'h1ACA;    //value='d 6858;             
          'd0918 : value = 'h1ACE;    //value='d 6862;             
          'd0919 : value = 'h1AD2;    //value='d 6866;             
          'd0920 : value = 'h1AD6;    //value='d 6870;             
          'd0921 : value = 'h1ADA;    //value='d 6874;             
          'd0922 : value = 'h1ADD;    //value='d 6877;             
          'd0923 : value = 'h1AE1;    //value='d 6881;             
          'd0924 : value = 'h1AE5;    //value='d 6885;             
          'd0925 : value = 'h1AE9;    //value='d 6889;             
          'd0926 : value = 'h1AED;    //value='d 6893;             
          'd0927 : value = 'h1AF1;    //value='d 6897;             
          'd0928 : value = 'h1AF5;    //value='d 6901;             
          'd0929 : value = 'h1AF9;    //value='d 6905;             
          'd0930 : value = 'h1AFC;    //value='d 6908;             
          'd0931 : value = 'h1B00;    //value='d 6912;             
          'd0932 : value = 'h1B04;    //value='d 6916;             
          'd0933 : value = 'h1B08;    //value='d 6920;             
          'd0934 : value = 'h1B0C;    //value='d 6924;             
          'd0935 : value = 'h1B10;    //value='d 6928;             
          'd0936 : value = 'h1B14;    //value='d 6932;             
          'd0937 : value = 'h1B18;    //value='d 6936;             
          'd0938 : value = 'h1B1C;    //value='d 6940;             
          'd0939 : value = 'h1B1F;    //value='d 6943;             
          'd0940 : value = 'h1B23;    //value='d 6947;             
          'd0941 : value = 'h1B27;    //value='d 6951;             
          'd0942 : value = 'h1B2B;    //value='d 6955;             
          'd0943 : value = 'h1B2F;    //value='d 6959;             
          'd0944 : value = 'h1B33;    //value='d 6963;             
          'd0945 : value = 'h1B37;    //value='d 6967;             
          'd0946 : value = 'h1B3B;    //value='d 6971;             
          'd0947 : value = 'h1B3F;    //value='d 6975;             
          'd0948 : value = 'h1B43;    //value='d 6979;             
          'd0949 : value = 'h1B47;    //value='d 6983;             
          'd0950 : value = 'h1B4B;    //value='d 6987;             
          'd0951 : value = 'h1B4E;    //value='d 6990;             
          'd0952 : value = 'h1B52;    //value='d 6994;             
          'd0953 : value = 'h1B56;    //value='d 6998;             
          'd0954 : value = 'h1B5A;    //value='d 7002;             
          'd0955 : value = 'h1B5E;    //value='d 7006;             
          'd0956 : value = 'h1B62;    //value='d 7010;             
          'd0957 : value = 'h1B66;    //value='d 7014;             
          'd0958 : value = 'h1B6A;    //value='d 7018;             
          'd0959 : value = 'h1B6E;    //value='d 7022;             
          'd0960 : value = 'h1B72;    //value='d 7026;             
          'd0961 : value = 'h1B76;    //value='d 7030;             
          'd0962 : value = 'h1B7A;    //value='d 7034;             
          'd0963 : value = 'h1B7E;    //value='d 7038;             
          'd0964 : value = 'h1B82;    //value='d 7042;             
          'd0965 : value = 'h1B86;    //value='d 7046;             
          'd0966 : value = 'h1B8A;    //value='d 7050;             
          'd0967 : value = 'h1B8E;    //value='d 7054;             
          'd0968 : value = 'h1B92;    //value='d 7058;             
          'd0969 : value = 'h1B96;    //value='d 7062;             
          'd0970 : value = 'h1B9A;    //value='d 7066;             
          'd0971 : value = 'h1B9E;    //value='d 7070;             
          'd0972 : value = 'h1BA1;    //value='d 7073;             
          'd0973 : value = 'h1BA5;    //value='d 7077;             
          'd0974 : value = 'h1BA9;    //value='d 7081;             
          'd0975 : value = 'h1BAD;    //value='d 7085;             
          'd0976 : value = 'h1BB1;    //value='d 7089;             
          'd0977 : value = 'h1BB5;    //value='d 7093;             
          'd0978 : value = 'h1BB9;    //value='d 7097;             
          'd0979 : value = 'h1BBD;    //value='d 7101;             
          'd0980 : value = 'h1BC1;    //value='d 7105;             
          'd0981 : value = 'h1BC5;    //value='d 7109;             
          'd0982 : value = 'h1BC9;    //value='d 7113;             
          'd0983 : value = 'h1BCD;    //value='d 7117;             
          'd0984 : value = 'h1BD1;    //value='d 7121;             
          'd0985 : value = 'h1BD5;    //value='d 7125;             
          'd0986 : value = 'h1BD9;    //value='d 7129;             
          'd0987 : value = 'h1BDD;    //value='d 7133;             
          'd0988 : value = 'h1BE1;    //value='d 7137;             
          'd0989 : value = 'h1BE5;    //value='d 7141;             
          'd0990 : value = 'h1BE9;    //value='d 7145;             
          'd0991 : value = 'h1BED;    //value='d 7149;             
          'd0992 : value = 'h1BF1;    //value='d 7153;             
          'd0993 : value = 'h1BF5;    //value='d 7157;             
          'd0994 : value = 'h1BFA;    //value='d 7162;             
          'd0995 : value = 'h1BFE;    //value='d 7166;             
          'd0996 : value = 'h1C02;    //value='d 7170;             
          'd0997 : value = 'h1C06;    //value='d 7174;             
          'd0998 : value = 'h1C0A;    //value='d 7178;             
          'd0999 : value = 'h1C0E;    //value='d 7182;             
          'd1000 : value = 'h1C12;    //value='d 7186;             
          'd1001 : value = 'h1C16;    //value='d 7190;             
          'd1002 : value = 'h1C1A;    //value='d 7194;             
          'd1003 : value = 'h1C1E;    //value='d 7198;             
          'd1004 : value = 'h1C22;    //value='d 7202;             
          'd1005 : value = 'h1C26;    //value='d 7206;             
          'd1006 : value = 'h1C2A;    //value='d 7210;             
          'd1007 : value = 'h1C2E;    //value='d 7214;             
          'd1008 : value = 'h1C32;    //value='d 7218;             
          'd1009 : value = 'h1C36;    //value='d 7222;             
          'd1010 : value = 'h1C3A;    //value='d 7226;             
          'd1011 : value = 'h1C3E;    //value='d 7230;             
          'd1012 : value = 'h1C42;    //value='d 7234;             
          'd1013 : value = 'h1C46;    //value='d 7238;             
          'd1014 : value = 'h1C4B;    //value='d 7243;             
          'd1015 : value = 'h1C4F;    //value='d 7247;             
          'd1016 : value = 'h1C53;    //value='d 7251;             
          'd1017 : value = 'h1C57;    //value='d 7255;             
          'd1018 : value = 'h1C5B;    //value='d 7259;             
          'd1019 : value = 'h1C5F;    //value='d 7263;             
          'd1020 : value = 'h1C63;    //value='d 7267;             
          'd1021 : value = 'h1C67;    //value='d 7271;             
          'd1022 : value = 'h1C6B;    //value='d 7275;             
          'd1023 : value = 'h1C6F;    //value='d 7279;             
          'd1024 : value = 'h1C73;    //value='d 7283;             
          'd1025 : value = 'h1C77;    //value='d 7287;             
          'd1026 : value = 'h1C7C;    //value='d 7292;             
          'd1027 : value = 'h1C80;    //value='d 7296;             
          'd1028 : value = 'h1C84;    //value='d 7300;             
          'd1029 : value = 'h1C88;    //value='d 7304;             
          'd1030 : value = 'h1C8C;    //value='d 7308;             
          'd1031 : value = 'h1C90;    //value='d 7312;             
          'd1032 : value = 'h1C94;    //value='d 7316;             
          'd1033 : value = 'h1C98;    //value='d 7320;             
          'd1034 : value = 'h1C9C;    //value='d 7324;             
          'd1035 : value = 'h1CA1;    //value='d 7329;             
          'd1036 : value = 'h1CA5;    //value='d 7333;             
          'd1037 : value = 'h1CA9;    //value='d 7337;             
          'd1038 : value = 'h1CAD;    //value='d 7341;             
          'd1039 : value = 'h1CB1;    //value='d 7345;             
          'd1040 : value = 'h1CB5;    //value='d 7349;             
          'd1041 : value = 'h1CB9;    //value='d 7353;             
          'd1042 : value = 'h1CBD;    //value='d 7357;             
          'd1043 : value = 'h1CC2;    //value='d 7362;             
          'd1044 : value = 'h1CC6;    //value='d 7366;             
          'd1045 : value = 'h1CCA;    //value='d 7370;             
          'd1046 : value = 'h1CCE;    //value='d 7374;             
          'd1047 : value = 'h1CD2;    //value='d 7378;             
          'd1048 : value = 'h1CD6;    //value='d 7382;             
          'd1049 : value = 'h1CDA;    //value='d 7386;             
          'd1050 : value = 'h1CDF;    //value='d 7391;             
          'd1051 : value = 'h1CE3;    //value='d 7395;             
          'd1052 : value = 'h1CE7;    //value='d 7399;             
          'd1053 : value = 'h1CEB;    //value='d 7403;             
          'd1054 : value = 'h1CEF;    //value='d 7407;             
          'd1055 : value = 'h1CF3;    //value='d 7411;             
          'd1056 : value = 'h1CF8;    //value='d 7416;             
          'd1057 : value = 'h1CFC;    //value='d 7420;             
          'd1058 : value = 'h1D00;    //value='d 7424;             
          'd1059 : value = 'h1D04;    //value='d 7428;             
          'd1060 : value = 'h1D08;    //value='d 7432;             
          'd1061 : value = 'h1D0C;    //value='d 7436;             
          'd1062 : value = 'h1D11;    //value='d 7441;             
          'd1063 : value = 'h1D15;    //value='d 7445;             
          'd1064 : value = 'h1D19;    //value='d 7449;             
          'd1065 : value = 'h1D1D;    //value='d 7453;             
          'd1066 : value = 'h1D21;    //value='d 7457;             
          'd1067 : value = 'h1D26;    //value='d 7462;             
          'd1068 : value = 'h1D2A;    //value='d 7466;             
          'd1069 : value = 'h1D2E;    //value='d 7470;             
          'd1070 : value = 'h1D32;    //value='d 7474;             
          'd1071 : value = 'h1D36;    //value='d 7478;             
          'd1072 : value = 'h1D3B;    //value='d 7483;             
          'd1073 : value = 'h1D3F;    //value='d 7487;             
          'd1074 : value = 'h1D43;    //value='d 7491;             
          'd1075 : value = 'h1D47;    //value='d 7495;             
          'd1076 : value = 'h1D4B;    //value='d 7499;             
          'd1077 : value = 'h1D50;    //value='d 7504;             
          'd1078 : value = 'h1D54;    //value='d 7508;             
          'd1079 : value = 'h1D58;    //value='d 7512;             
          'd1080 : value = 'h1D5C;    //value='d 7516;             
          'd1081 : value = 'h1D61;    //value='d 7521;             
          'd1082 : value = 'h1D65;    //value='d 7525;             
          'd1083 : value = 'h1D69;    //value='d 7529;             
          'd1084 : value = 'h1D6D;    //value='d 7533;             
          'd1085 : value = 'h1D71;    //value='d 7537;             
          'd1086 : value = 'h1D76;    //value='d 7542;             
          'd1087 : value = 'h1D7A;    //value='d 7546;             
          'd1088 : value = 'h1D7E;    //value='d 7550;             
          'd1089 : value = 'h1D82;    //value='d 7554;             
          'd1090 : value = 'h1D87;    //value='d 7559;             
          'd1091 : value = 'h1D8B;    //value='d 7563;             
          'd1092 : value = 'h1D8F;    //value='d 7567;             
          'd1093 : value = 'h1D93;    //value='d 7571;             
          'd1094 : value = 'h1D98;    //value='d 7576;             
          'd1095 : value = 'h1D9C;    //value='d 7580;             
          'd1096 : value = 'h1DA0;    //value='d 7584;             
          'd1097 : value = 'h1DA4;    //value='d 7588;             
          'd1098 : value = 'h1DA9;    //value='d 7593;             
          'd1099 : value = 'h1DAD;    //value='d 7597;             
          'd1100 : value = 'h1DB1;    //value='d 7601;             
          'd1101 : value = 'h1DB6;    //value='d 7606;             
          'd1102 : value = 'h1DBA;    //value='d 7610;             
          'd1103 : value = 'h1DBE;    //value='d 7614;             
          'd1104 : value = 'h1DC2;    //value='d 7618;             
          'd1105 : value = 'h1DC7;    //value='d 7623;             
          'd1106 : value = 'h1DCB;    //value='d 7627;             
          'd1107 : value = 'h1DCF;    //value='d 7631;             
          'd1108 : value = 'h1DD4;    //value='d 7636;             
          'd1109 : value = 'h1DD8;    //value='d 7640;             
          'd1110 : value = 'h1DDC;    //value='d 7644;             
          'd1111 : value = 'h1DE0;    //value='d 7648;             
          'd1112 : value = 'h1DE5;    //value='d 7653;             
          'd1113 : value = 'h1DE9;    //value='d 7657;             
          'd1114 : value = 'h1DED;    //value='d 7661;             
          'd1115 : value = 'h1DF2;    //value='d 7666;             
          'd1116 : value = 'h1DF6;    //value='d 7670;             
          'd1117 : value = 'h1DFA;    //value='d 7674;             
          'd1118 : value = 'h1DFF;    //value='d 7679;             
          'd1119 : value = 'h1E03;    //value='d 7683;             
          'd1120 : value = 'h1E07;    //value='d 7687;             
          'd1121 : value = 'h1E0C;    //value='d 7692;             
          'd1122 : value = 'h1E10;    //value='d 7696;             
          'd1123 : value = 'h1E14;    //value='d 7700;             
          'd1124 : value = 'h1E19;    //value='d 7705;             
          'd1125 : value = 'h1E1D;    //value='d 7709;             
          'd1126 : value = 'h1E21;    //value='d 7713;             
          'd1127 : value = 'h1E26;    //value='d 7718;             
          'd1128 : value = 'h1E2A;    //value='d 7722;             
          'd1129 : value = 'h1E2E;    //value='d 7726;             
          'd1130 : value = 'h1E33;    //value='d 7731;             
          'd1131 : value = 'h1E37;    //value='d 7735;             
          'd1132 : value = 'h1E3B;    //value='d 7739;             
          'd1133 : value = 'h1E40;    //value='d 7744;             
          'd1134 : value = 'h1E44;    //value='d 7748;             
          'd1135 : value = 'h1E48;    //value='d 7752;             
          'd1136 : value = 'h1E4D;    //value='d 7757;             
          'd1137 : value = 'h1E51;    //value='d 7761;             
          'd1138 : value = 'h1E55;    //value='d 7765;             
          'd1139 : value = 'h1E5A;    //value='d 7770;             
          'd1140 : value = 'h1E5E;    //value='d 7774;             
          'd1141 : value = 'h1E63;    //value='d 7779;             
          'd1142 : value = 'h1E67;    //value='d 7783;             
          'd1143 : value = 'h1E6B;    //value='d 7787;             
          'd1144 : value = 'h1E70;    //value='d 7792;             
          'd1145 : value = 'h1E74;    //value='d 7796;             
          'd1146 : value = 'h1E78;    //value='d 7800;             
          'd1147 : value = 'h1E7D;    //value='d 7805;             
          'd1148 : value = 'h1E81;    //value='d 7809;             
          'd1149 : value = 'h1E86;    //value='d 7814;             
          'd1150 : value = 'h1E8A;    //value='d 7818;             
          'd1151 : value = 'h1E8E;    //value='d 7822;             
          'd1152 : value = 'h1E93;    //value='d 7827;             
          'd1153 : value = 'h1E97;    //value='d 7831;             
          'd1154 : value = 'h1E9C;    //value='d 7836;             
          'd1155 : value = 'h1EA0;    //value='d 7840;             
          'd1156 : value = 'h1EA4;    //value='d 7844;             
          'd1157 : value = 'h1EA9;    //value='d 7849;             
          'd1158 : value = 'h1EAD;    //value='d 7853;             
          'd1159 : value = 'h1EB2;    //value='d 7858;             
          'd1160 : value = 'h1EB6;    //value='d 7862;             
          'd1161 : value = 'h1EBA;    //value='d 7866;             
          'd1162 : value = 'h1EBF;    //value='d 7871;             
          'd1163 : value = 'h1EC3;    //value='d 7875;             
          'd1164 : value = 'h1EC8;    //value='d 7880;             
          'd1165 : value = 'h1ECC;    //value='d 7884;             
          'd1166 : value = 'h1ED1;    //value='d 7889;             
          'd1167 : value = 'h1ED5;    //value='d 7893;             
          'd1168 : value = 'h1ED9;    //value='d 7897;             
          'd1169 : value = 'h1EDE;    //value='d 7902;             
          'd1170 : value = 'h1EE2;    //value='d 7906;             
          'd1171 : value = 'h1EE7;    //value='d 7911;             
          'd1172 : value = 'h1EEB;    //value='d 7915;             
          'd1173 : value = 'h1EF0;    //value='d 7920;             
          'd1174 : value = 'h1EF4;    //value='d 7924;             
          'd1175 : value = 'h1EF9;    //value='d 7929;             
          'd1176 : value = 'h1EFD;    //value='d 7933;             
          'd1177 : value = 'h1F02;    //value='d 7938;             
          'd1178 : value = 'h1F06;    //value='d 7942;             
          'd1179 : value = 'h1F0A;    //value='d 7946;             
          'd1180 : value = 'h1F0F;    //value='d 7951;             
          'd1181 : value = 'h1F13;    //value='d 7955;             
          'd1182 : value = 'h1F18;    //value='d 7960;             
          'd1183 : value = 'h1F1C;    //value='d 7964;             
          'd1184 : value = 'h1F21;    //value='d 7969;             
          'd1185 : value = 'h1F25;    //value='d 7973;             
          'd1186 : value = 'h1F2A;    //value='d 7978;             
          'd1187 : value = 'h1F2E;    //value='d 7982;             
          'd1188 : value = 'h1F33;    //value='d 7987;             
          'd1189 : value = 'h1F37;    //value='d 7991;             
          'd1190 : value = 'h1F3C;    //value='d 7996;             
          'd1191 : value = 'h1F40;    //value='d 8000;             
          'd1192 : value = 'h1F45;    //value='d 8005;             
          'd1193 : value = 'h1F49;    //value='d 8009;             
          'd1194 : value = 'h1F4E;    //value='d 8014;             
          'd1195 : value = 'h1F52;    //value='d 8018;             
          'd1196 : value = 'h1F57;    //value='d 8023;             
          'd1197 : value = 'h1F5B;    //value='d 8027;             
          'd1198 : value = 'h1F60;    //value='d 8032;             
          'd1199 : value = 'h1F64;    //value='d 8036;             
          'd1200 : value = 'h1F69;    //value='d 8041;             
          'd1201 : value = 'h1F6D;    //value='d 8045;             
          'd1202 : value = 'h1F72;    //value='d 8050;             
          'd1203 : value = 'h1F76;    //value='d 8054;             
          'd1204 : value = 'h1F7B;    //value='d 8059;             
          'd1205 : value = 'h1F7F;    //value='d 8063;             
          'd1206 : value = 'h1F84;    //value='d 8068;             
          'd1207 : value = 'h1F89;    //value='d 8073;             
          'd1208 : value = 'h1F8D;    //value='d 8077;             
          'd1209 : value = 'h1F92;    //value='d 8082;             
          'd1210 : value = 'h1F96;    //value='d 8086;             
          'd1211 : value = 'h1F9B;    //value='d 8091;             
          'd1212 : value = 'h1F9F;    //value='d 8095;             
          'd1213 : value = 'h1FA4;    //value='d 8100;             
          'd1214 : value = 'h1FA8;    //value='d 8104;             
          'd1215 : value = 'h1FAD;    //value='d 8109;             
          'd1216 : value = 'h1FB1;    //value='d 8113;             
          'd1217 : value = 'h1FB6;    //value='d 8118;             
          'd1218 : value = 'h1FBB;    //value='d 8123;             
          'd1219 : value = 'h1FBF;    //value='d 8127;             
          'd1220 : value = 'h1FC4;    //value='d 8132;             
          'd1221 : value = 'h1FC8;    //value='d 8136;             
          'd1222 : value = 'h1FCD;    //value='d 8141;             
          'd1223 : value = 'h1FD1;    //value='d 8145;             
          'd1224 : value = 'h1FD6;    //value='d 8150;             
          'd1225 : value = 'h1FDB;    //value='d 8155;             
          'd1226 : value = 'h1FDF;    //value='d 8159;             
          'd1227 : value = 'h1FE4;    //value='d 8164;             
          'd1228 : value = 'h1FE8;    //value='d 8168;             
          'd1229 : value = 'h1FED;    //value='d 8173;             
          'd1230 : value = 'h1FF2;    //value='d 8178;             
          'd1231 : value = 'h1FF6;    //value='d 8182;             
          'd1232 : value = 'h1FFB;    //value='d 8187;             
          'd1233 : value = 'h1FFF;    //value='d 8191;             
          'd1234 : value = 'h2004;    //value='d 8196;             
          'd1235 : value = 'h2009;    //value='d 8201;             
          'd1236 : value = 'h200D;    //value='d 8205;             
          'd1237 : value = 'h2012;    //value='d 8210;             
          'd1238 : value = 'h2016;    //value='d 8214;             
          'd1239 : value = 'h201B;    //value='d 8219;             
          'd1240 : value = 'h2020;    //value='d 8224;             
          'd1241 : value = 'h2024;    //value='d 8228;             
          'd1242 : value = 'h2029;    //value='d 8233;             
          'd1243 : value = 'h202E;    //value='d 8238;             
          'd1244 : value = 'h2032;    //value='d 8242;             
          'd1245 : value = 'h2037;    //value='d 8247;             
          'd1246 : value = 'h203B;    //value='d 8251;             
          'd1247 : value = 'h2040;    //value='d 8256;             
          'd1248 : value = 'h2045;    //value='d 8261;             
          'd1249 : value = 'h2049;    //value='d 8265;             
          'd1250 : value = 'h204E;    //value='d 8270;             
          'd1251 : value = 'h2053;    //value='d 8275;             
          'd1252 : value = 'h2057;    //value='d 8279;             
          'd1253 : value = 'h205C;    //value='d 8284;             
          'd1254 : value = 'h2061;    //value='d 8289;             
          'd1255 : value = 'h2065;    //value='d 8293;             
          'd1256 : value = 'h206A;    //value='d 8298;             
          'd1257 : value = 'h206F;    //value='d 8303;             
          'd1258 : value = 'h2073;    //value='d 8307;             
          'd1259 : value = 'h2078;    //value='d 8312;             
          'd1260 : value = 'h207D;    //value='d 8317;             
          'd1261 : value = 'h2081;    //value='d 8321;             
          'd1262 : value = 'h2086;    //value='d 8326;             
          'd1263 : value = 'h208B;    //value='d 8331;             
          'd1264 : value = 'h208F;    //value='d 8335;             
          'd1265 : value = 'h2094;    //value='d 8340;             
          'd1266 : value = 'h2099;    //value='d 8345;             
          'd1267 : value = 'h209D;    //value='d 8349;             
          'd1268 : value = 'h20A2;    //value='d 8354;             
          'd1269 : value = 'h20A7;    //value='d 8359;             
          'd1270 : value = 'h20AC;    //value='d 8364;             
          'd1271 : value = 'h20B0;    //value='d 8368;             
          'd1272 : value = 'h20B5;    //value='d 8373;             
          'd1273 : value = 'h20BA;    //value='d 8378;             
          'd1274 : value = 'h20BE;    //value='d 8382;             
          'd1275 : value = 'h20C3;    //value='d 8387;             
          'd1276 : value = 'h20C8;    //value='d 8392;             
          'd1277 : value = 'h20CD;    //value='d 8397;             
          'd1278 : value = 'h20D1;    //value='d 8401;             
          'd1279 : value = 'h20D6;    //value='d 8406;             
          'd1280 : value = 'h20DB;    //value='d 8411;             
          'd1281 : value = 'h20DF;    //value='d 8415;             
          'd1282 : value = 'h20E4;    //value='d 8420;             
          'd1283 : value = 'h20E9;    //value='d 8425;             
          'd1284 : value = 'h20EE;    //value='d 8430;             
          'd1285 : value = 'h20F2;    //value='d 8434;             
          'd1286 : value = 'h20F7;    //value='d 8439;             
          'd1287 : value = 'h20FC;    //value='d 8444;             
          'd1288 : value = 'h2101;    //value='d 8449;             
          'd1289 : value = 'h2105;    //value='d 8453;             
          'd1290 : value = 'h210A;    //value='d 8458;             
          'd1291 : value = 'h210F;    //value='d 8463;             
          'd1292 : value = 'h2114;    //value='d 8468;             
          'd1293 : value = 'h2118;    //value='d 8472;             
          'd1294 : value = 'h211D;    //value='d 8477;             
          'd1295 : value = 'h2122;    //value='d 8482;             
          'd1296 : value = 'h2127;    //value='d 8487;             
          'd1297 : value = 'h212C;    //value='d 8492;             
          'd1298 : value = 'h2130;    //value='d 8496;             
          'd1299 : value = 'h2135;    //value='d 8501;             
          'd1300 : value = 'h213A;    //value='d 8506;             
          'd1301 : value = 'h213F;    //value='d 8511;             
          'd1302 : value = 'h2143;    //value='d 8515;             
          'd1303 : value = 'h2148;    //value='d 8520;             
          'd1304 : value = 'h214D;    //value='d 8525;             
          'd1305 : value = 'h2152;    //value='d 8530;             
          'd1306 : value = 'h2157;    //value='d 8535;             
          'd1307 : value = 'h215B;    //value='d 8539;             
          'd1308 : value = 'h2160;    //value='d 8544;             
          'd1309 : value = 'h2165;    //value='d 8549;             
          'd1310 : value = 'h216A;    //value='d 8554;             
          'd1311 : value = 'h216F;    //value='d 8559;             
          'd1312 : value = 'h2173;    //value='d 8563;             
          'd1313 : value = 'h2178;    //value='d 8568;             
          'd1314 : value = 'h217D;    //value='d 8573;             
          'd1315 : value = 'h2182;    //value='d 8578;             
          'd1316 : value = 'h2187;    //value='d 8583;             
          'd1317 : value = 'h218C;    //value='d 8588;             
          'd1318 : value = 'h2190;    //value='d 8592;             
          'd1319 : value = 'h2195;    //value='d 8597;             
          'd1320 : value = 'h219A;    //value='d 8602;             
          'd1321 : value = 'h219F;    //value='d 8607;             
          'd1322 : value = 'h21A4;    //value='d 8612;             
          'd1323 : value = 'h21A9;    //value='d 8617;             
          'd1324 : value = 'h21AD;    //value='d 8621;             
          'd1325 : value = 'h21B2;    //value='d 8626;             
          'd1326 : value = 'h21B7;    //value='d 8631;             
          'd1327 : value = 'h21BC;    //value='d 8636;             
          'd1328 : value = 'h21C1;    //value='d 8641;             
          'd1329 : value = 'h21C6;    //value='d 8646;             
          'd1330 : value = 'h21CB;    //value='d 8651;             
          'd1331 : value = 'h21CF;    //value='d 8655;             
          'd1332 : value = 'h21D4;    //value='d 8660;             
          'd1333 : value = 'h21D9;    //value='d 8665;             
          'd1334 : value = 'h21DE;    //value='d 8670;             
          'd1335 : value = 'h21E3;    //value='d 8675;             
          'd1336 : value = 'h21E8;    //value='d 8680;             
          'd1337 : value = 'h21ED;    //value='d 8685;             
          'd1338 : value = 'h21F2;    //value='d 8690;             
          'd1339 : value = 'h21F6;    //value='d 8694;             
          'd1340 : value = 'h21FB;    //value='d 8699;             
          'd1341 : value = 'h2200;    //value='d 8704;             
          'd1342 : value = 'h2205;    //value='d 8709;             
          'd1343 : value = 'h220A;    //value='d 8714;             
          'd1344 : value = 'h220F;    //value='d 8719;             
          'd1345 : value = 'h2214;    //value='d 8724;             
          'd1346 : value = 'h2219;    //value='d 8729;             
          'd1347 : value = 'h221E;    //value='d 8734;             
          'd1348 : value = 'h2222;    //value='d 8738;             
          'd1349 : value = 'h2227;    //value='d 8743;             
          'd1350 : value = 'h222C;    //value='d 8748;             
          'd1351 : value = 'h2231;    //value='d 8753;             
          'd1352 : value = 'h2236;    //value='d 8758;             
          'd1353 : value = 'h223B;    //value='d 8763;             
          'd1354 : value = 'h2240;    //value='d 8768;             
          'd1355 : value = 'h2245;    //value='d 8773;             
          'd1356 : value = 'h224A;    //value='d 8778;             
          'd1357 : value = 'h224F;    //value='d 8783;             
          'd1358 : value = 'h2254;    //value='d 8788;             
          'd1359 : value = 'h2259;    //value='d 8793;             
          'd1360 : value = 'h225E;    //value='d 8798;             
          'd1361 : value = 'h2263;    //value='d 8803;             
          'd1362 : value = 'h2268;    //value='d 8808;             
          'd1363 : value = 'h226C;    //value='d 8812;             
          'd1364 : value = 'h2271;    //value='d 8817;             
          'd1365 : value = 'h2276;    //value='d 8822;             
          'd1366 : value = 'h227B;    //value='d 8827;             
          'd1367 : value = 'h2280;    //value='d 8832;             
          'd1368 : value = 'h2285;    //value='d 8837;             
          'd1369 : value = 'h228A;    //value='d 8842;             
          'd1370 : value = 'h228F;    //value='d 8847;             
          'd1371 : value = 'h2294;    //value='d 8852;             
          'd1372 : value = 'h2299;    //value='d 8857;             
          'd1373 : value = 'h229E;    //value='d 8862;             
          'd1374 : value = 'h22A3;    //value='d 8867;             
          'd1375 : value = 'h22A8;    //value='d 8872;             
          'd1376 : value = 'h22AD;    //value='d 8877;             
          'd1377 : value = 'h22B2;    //value='d 8882;             
          'd1378 : value = 'h22B7;    //value='d 8887;             
          'd1379 : value = 'h22BC;    //value='d 8892;             
          'd1380 : value = 'h22C1;    //value='d 8897;             
          'd1381 : value = 'h22C6;    //value='d 8902;             
          'd1382 : value = 'h22CB;    //value='d 8907;             
          'd1383 : value = 'h22D0;    //value='d 8912;             
          'd1384 : value = 'h22D5;    //value='d 8917;             
          'd1385 : value = 'h22DA;    //value='d 8922;             
          'd1386 : value = 'h22DF;    //value='d 8927;             
          'd1387 : value = 'h22E4;    //value='d 8932;             
          'd1388 : value = 'h22E9;    //value='d 8937;             
          'd1389 : value = 'h22EE;    //value='d 8942;             
          'd1390 : value = 'h22F3;    //value='d 8947;             
          'd1391 : value = 'h22F8;    //value='d 8952;             
          'd1392 : value = 'h22FD;    //value='d 8957;             
          'd1393 : value = 'h2302;    //value='d 8962;             
          'd1394 : value = 'h2307;    //value='d 8967;             
          'd1395 : value = 'h230C;    //value='d 8972;             
          'd1396 : value = 'h2312;    //value='d 8978;             
          'd1397 : value = 'h2317;    //value='d 8983;             
          'd1398 : value = 'h231C;    //value='d 8988;             
          'd1399 : value = 'h2321;    //value='d 8993;             
          'd1400 : value = 'h2326;    //value='d 8998;             
          'd1401 : value = 'h232B;    //value='d 9003;             
          'd1402 : value = 'h2330;    //value='d 9008;             
          'd1403 : value = 'h2335;    //value='d 9013;             
          'd1404 : value = 'h233A;    //value='d 9018;             
          'd1405 : value = 'h233F;    //value='d 9023;             
          'd1406 : value = 'h2344;    //value='d 9028;             
          'd1407 : value = 'h2349;    //value='d 9033;             
          'd1408 : value = 'h234E;    //value='d 9038;             
          'd1409 : value = 'h2353;    //value='d 9043;             
          'd1410 : value = 'h2358;    //value='d 9048;             
          'd1411 : value = 'h235E;    //value='d 9054;             
          'd1412 : value = 'h2363;    //value='d 9059;             
          'd1413 : value = 'h2368;    //value='d 9064;             
          'd1414 : value = 'h236D;    //value='d 9069;             
          'd1415 : value = 'h2372;    //value='d 9074;             
          'd1416 : value = 'h2377;    //value='d 9079;             
          'd1417 : value = 'h237C;    //value='d 9084;             
          'd1418 : value = 'h2381;    //value='d 9089;             
          'd1419 : value = 'h2386;    //value='d 9094;             
          'd1420 : value = 'h238B;    //value='d 9099;             
          'd1421 : value = 'h2391;    //value='d 9105;             
          'd1422 : value = 'h2396;    //value='d 9110;             
          'd1423 : value = 'h239B;    //value='d 9115;             
          'd1424 : value = 'h23A0;    //value='d 9120;             
          'd1425 : value = 'h23A5;    //value='d 9125;             
          'd1426 : value = 'h23AA;    //value='d 9130;             
          'd1427 : value = 'h23AF;    //value='d 9135;             
          'd1428 : value = 'h23B4;    //value='d 9140;             
          'd1429 : value = 'h23BA;    //value='d 9146;             
          'd1430 : value = 'h23BF;    //value='d 9151;             
          'd1431 : value = 'h23C4;    //value='d 9156;             
          'd1432 : value = 'h23C9;    //value='d 9161;             
          'd1433 : value = 'h23CE;    //value='d 9166;             
          'd1434 : value = 'h23D3;    //value='d 9171;             
          'd1435 : value = 'h23D9;    //value='d 9177;             
          'd1436 : value = 'h23DE;    //value='d 9182;             
          'd1437 : value = 'h23E3;    //value='d 9187;             
          'd1438 : value = 'h23E8;    //value='d 9192;             
          'd1439 : value = 'h23ED;    //value='d 9197;             
          'd1440 : value = 'h23F2;    //value='d 9202;             
          'd1441 : value = 'h23F8;    //value='d 9208;             
          'd1442 : value = 'h23FD;    //value='d 9213;             
          'd1443 : value = 'h2402;    //value='d 9218;             
          'd1444 : value = 'h2407;    //value='d 9223;             
          'd1445 : value = 'h240C;    //value='d 9228;             
          'd1446 : value = 'h2411;    //value='d 9233;             
          'd1447 : value = 'h2417;    //value='d 9239;             
          'd1448 : value = 'h241C;    //value='d 9244;             
          'd1449 : value = 'h2421;    //value='d 9249;             
          'd1450 : value = 'h2426;    //value='d 9254;             
          'd1451 : value = 'h242B;    //value='d 9259;             
          'd1452 : value = 'h2431;    //value='d 9265;             
          'd1453 : value = 'h2436;    //value='d 9270;             
          'd1454 : value = 'h243B;    //value='d 9275;             
          'd1455 : value = 'h2440;    //value='d 9280;             
          'd1456 : value = 'h2446;    //value='d 9286;             
          'd1457 : value = 'h244B;    //value='d 9291;             
          'd1458 : value = 'h2450;    //value='d 9296;             
          'd1459 : value = 'h2455;    //value='d 9301;             
          'd1460 : value = 'h245A;    //value='d 9306;             
          'd1461 : value = 'h2460;    //value='d 9312;             
          'd1462 : value = 'h2465;    //value='d 9317;             
          'd1463 : value = 'h246A;    //value='d 9322;             
          'd1464 : value = 'h246F;    //value='d 9327;             
          'd1465 : value = 'h2475;    //value='d 9333;             
          'd1466 : value = 'h247A;    //value='d 9338;             
          'd1467 : value = 'h247F;    //value='d 9343;             
          'd1468 : value = 'h2484;    //value='d 9348;             
          'd1469 : value = 'h248A;    //value='d 9354;             
          'd1470 : value = 'h248F;    //value='d 9359;             
          'd1471 : value = 'h2494;    //value='d 9364;             
          'd1472 : value = 'h2499;    //value='d 9369;             
          'd1473 : value = 'h249F;    //value='d 9375;             
          'd1474 : value = 'h24A4;    //value='d 9380;             
          'd1475 : value = 'h24A9;    //value='d 9385;             
          'd1476 : value = 'h24AE;    //value='d 9390;             
          'd1477 : value = 'h24B4;    //value='d 9396;             
          'd1478 : value = 'h24B9;    //value='d 9401;             
          'd1479 : value = 'h24BE;    //value='d 9406;             
          'd1480 : value = 'h24C4;    //value='d 9412;             
          'd1481 : value = 'h24C9;    //value='d 9417;             
          'd1482 : value = 'h24CE;    //value='d 9422;             
          'd1483 : value = 'h24D4;    //value='d 9428;             
          'd1484 : value = 'h24D9;    //value='d 9433;             
          'd1485 : value = 'h24DE;    //value='d 9438;             
          'd1486 : value = 'h24E3;    //value='d 9443;             
          'd1487 : value = 'h24E9;    //value='d 9449;             
          'd1488 : value = 'h24EE;    //value='d 9454;             
          'd1489 : value = 'h24F3;    //value='d 9459;             
          'd1490 : value = 'h24F9;    //value='d 9465;             
          'd1491 : value = 'h24FE;    //value='d 9470;             
          'd1492 : value = 'h2503;    //value='d 9475;             
          'd1493 : value = 'h2509;    //value='d 9481;             
          'd1494 : value = 'h250E;    //value='d 9486;             
          'd1495 : value = 'h2513;    //value='d 9491;             
          'd1496 : value = 'h2519;    //value='d 9497;             
          'd1497 : value = 'h251E;    //value='d 9502;             
          'd1498 : value = 'h2523;    //value='d 9507;             
          'd1499 : value = 'h2529;    //value='d 9513;             
          'd1500 : value = 'h252E;    //value='d 9518;             
          'd1501 : value = 'h2533;    //value='d 9523;             
          'd1502 : value = 'h2539;    //value='d 9529;             
          'd1503 : value = 'h253E;    //value='d 9534;             
          'd1504 : value = 'h2543;    //value='d 9539;             
          'd1505 : value = 'h2549;    //value='d 9545;             
          'd1506 : value = 'h254E;    //value='d 9550;             
          'd1507 : value = 'h2554;    //value='d 9556;             
          'd1508 : value = 'h2559;    //value='d 9561;             
          'd1509 : value = 'h255E;    //value='d 9566;             
          'd1510 : value = 'h2564;    //value='d 9572;             
          'd1511 : value = 'h2569;    //value='d 9577;             
          'd1512 : value = 'h256E;    //value='d 9582;             
          'd1513 : value = 'h2574;    //value='d 9588;             
          'd1514 : value = 'h2579;    //value='d 9593;             
          'd1515 : value = 'h257F;    //value='d 9599;             
          'd1516 : value = 'h2584;    //value='d 9604;             
          'd1517 : value = 'h2589;    //value='d 9609;             
          'd1518 : value = 'h258F;    //value='d 9615;             
          'd1519 : value = 'h2594;    //value='d 9620;             
          'd1520 : value = 'h259A;    //value='d 9626;             
          'd1521 : value = 'h259F;    //value='d 9631;             
          'd1522 : value = 'h25A5;    //value='d 9637;             
          'd1523 : value = 'h25AA;    //value='d 9642;             
          'd1524 : value = 'h25AF;    //value='d 9647;             
          'd1525 : value = 'h25B5;    //value='d 9653;             
          'd1526 : value = 'h25BA;    //value='d 9658;             
          'd1527 : value = 'h25C0;    //value='d 9664;             
          'd1528 : value = 'h25C5;    //value='d 9669;             
          'd1529 : value = 'h25CA;    //value='d 9674;             
          'd1530 : value = 'h25D0;    //value='d 9680;             
          'd1531 : value = 'h25D5;    //value='d 9685;             
          'd1532 : value = 'h25DB;    //value='d 9691;             
          'd1533 : value = 'h25E0;    //value='d 9696;             
          'd1534 : value = 'h25E6;    //value='d 9702;             
          'd1535 : value = 'h25EB;    //value='d 9707;             
          'd1536 : value = 'h25F1;    //value='d 9713;             
          'd1537 : value = 'h25F6;    //value='d 9718;             
          'd1538 : value = 'h25FC;    //value='d 9724;             
          'd1539 : value = 'h2601;    //value='d 9729;             
          'd1540 : value = 'h2607;    //value='d 9735;             
          'd1541 : value = 'h260C;    //value='d 9740;             
          'd1542 : value = 'h2611;    //value='d 9745;             
          'd1543 : value = 'h2617;    //value='d 9751;             
          'd1544 : value = 'h261C;    //value='d 9756;             
          'd1545 : value = 'h2622;    //value='d 9762;             
          'd1546 : value = 'h2627;    //value='d 9767;             
          'd1547 : value = 'h262D;    //value='d 9773;             
          'd1548 : value = 'h2632;    //value='d 9778;             
          'd1549 : value = 'h2638;    //value='d 9784;             
          'd1550 : value = 'h263D;    //value='d 9789;             
          'd1551 : value = 'h2643;    //value='d 9795;             
          'd1552 : value = 'h2648;    //value='d 9800;             
          'd1553 : value = 'h264E;    //value='d 9806;             
          'd1554 : value = 'h2653;    //value='d 9811;             
          'd1555 : value = 'h2659;    //value='d 9817;             
          'd1556 : value = 'h265E;    //value='d 9822;             
          'd1557 : value = 'h2664;    //value='d 9828;             
          'd1558 : value = 'h266A;    //value='d 9834;             
          'd1559 : value = 'h266F;    //value='d 9839;             
          'd1560 : value = 'h2675;    //value='d 9845;             
          'd1561 : value = 'h267A;    //value='d 9850;             
          'd1562 : value = 'h2680;    //value='d 9856;             
          'd1563 : value = 'h2685;    //value='d 9861;             
          'd1564 : value = 'h268B;    //value='d 9867;             
          'd1565 : value = 'h2690;    //value='d 9872;             
          'd1566 : value = 'h2696;    //value='d 9878;             
          'd1567 : value = 'h269B;    //value='d 9883;             
          'd1568 : value = 'h26A1;    //value='d 9889;             
          'd1569 : value = 'h26A7;    //value='d 9895;             
          'd1570 : value = 'h26AC;    //value='d 9900;             
          'd1571 : value = 'h26B2;    //value='d 9906;             
          'd1572 : value = 'h26B7;    //value='d 9911;             
          'd1573 : value = 'h26BD;    //value='d 9917;             
          'd1574 : value = 'h26C2;    //value='d 9922;             
          'd1575 : value = 'h26C8;    //value='d 9928;             
          'd1576 : value = 'h26CE;    //value='d 9934;             
          'd1577 : value = 'h26D3;    //value='d 9939;             
          'd1578 : value = 'h26D9;    //value='d 9945;             
          'd1579 : value = 'h26DE;    //value='d 9950;             
          'd1580 : value = 'h26E4;    //value='d 9956;             
          'd1581 : value = 'h26E9;    //value='d 9961;             
          'd1582 : value = 'h26EF;    //value='d 9967;             
          'd1583 : value = 'h26F5;    //value='d 9973;             
          'd1584 : value = 'h26FA;    //value='d 9978;             
          'd1585 : value = 'h2700;    //value='d 9984;             
          'd1586 : value = 'h2706;    //value='d 9990;             
          'd1587 : value = 'h270B;    //value='d 9995;             
          'd1588 : value = 'h2711;    //value='d10001;             
          'd1589 : value = 'h2716;    //value='d10006;             
          'd1590 : value = 'h271C;    //value='d10012;             
          'd1591 : value = 'h2722;    //value='d10018;             
          'd1592 : value = 'h2727;    //value='d10023;             
          'd1593 : value = 'h272D;    //value='d10029;             
          'd1594 : value = 'h2733;    //value='d10035;             
          'd1595 : value = 'h2738;    //value='d10040;             
          'd1596 : value = 'h273E;    //value='d10046;             
          'd1597 : value = 'h2744;    //value='d10052;             
          'd1598 : value = 'h2749;    //value='d10057;             
          'd1599 : value = 'h274F;    //value='d10063;             
          'd1600 : value = 'h2754;    //value='d10068;             
          'd1601 : value = 'h275A;    //value='d10074;             
          'd1602 : value = 'h2760;    //value='d10080;             
          'd1603 : value = 'h2765;    //value='d10085;             
          'd1604 : value = 'h276B;    //value='d10091;             
          'd1605 : value = 'h2771;    //value='d10097;             
          'd1606 : value = 'h2776;    //value='d10102;             
          'd1607 : value = 'h277C;    //value='d10108;             
          'd1608 : value = 'h2782;    //value='d10114;             
          'd1609 : value = 'h2788;    //value='d10120;             
          'd1610 : value = 'h278D;    //value='d10125;             
          'd1611 : value = 'h2793;    //value='d10131;             
          'd1612 : value = 'h2799;    //value='d10137;             
          'd1613 : value = 'h279E;    //value='d10142;             
          'd1614 : value = 'h27A4;    //value='d10148;             
          'd1615 : value = 'h27AA;    //value='d10154;             
          'd1616 : value = 'h27AF;    //value='d10159;             
          'd1617 : value = 'h27B5;    //value='d10165;             
          'd1618 : value = 'h27BB;    //value='d10171;             
          'd1619 : value = 'h27C1;    //value='d10177;             
          'd1620 : value = 'h27C6;    //value='d10182;             
          'd1621 : value = 'h27CC;    //value='d10188;             
          'd1622 : value = 'h27D2;    //value='d10194;             
          'd1623 : value = 'h27D8;    //value='d10200;             
          'd1624 : value = 'h27DD;    //value='d10205;             
          'd1625 : value = 'h27E3;    //value='d10211;             
          'd1626 : value = 'h27E9;    //value='d10217;             
          'd1627 : value = 'h27EE;    //value='d10222;             
          'd1628 : value = 'h27F4;    //value='d10228;             
          'd1629 : value = 'h27FA;    //value='d10234;             
          'd1630 : value = 'h2800;    //value='d10240;             
          'd1631 : value = 'h2805;    //value='d10245;             
          'd1632 : value = 'h280B;    //value='d10251;             
          'd1633 : value = 'h2811;    //value='d10257;             
          'd1634 : value = 'h2817;    //value='d10263;             
          'd1635 : value = 'h281D;    //value='d10269;             
          'd1636 : value = 'h2822;    //value='d10274;             
          'd1637 : value = 'h2828;    //value='d10280;             
          'd1638 : value = 'h282E;    //value='d10286;             
          'd1639 : value = 'h2834;    //value='d10292;             
          'd1640 : value = 'h2839;    //value='d10297;             
          'd1641 : value = 'h283F;    //value='d10303;             
          'd1642 : value = 'h2845;    //value='d10309;             
          'd1643 : value = 'h284B;    //value='d10315;             
          'd1644 : value = 'h2851;    //value='d10321;             
          'd1645 : value = 'h2856;    //value='d10326;             
          'd1646 : value = 'h285C;    //value='d10332;             
          'd1647 : value = 'h2862;    //value='d10338;             
          'd1648 : value = 'h2868;    //value='d10344;             
          'd1649 : value = 'h286E;    //value='d10350;             
          'd1650 : value = 'h2873;    //value='d10355;             
          'd1651 : value = 'h2879;    //value='d10361;             
          'd1652 : value = 'h287F;    //value='d10367;             
          'd1653 : value = 'h2885;    //value='d10373;             
          'd1654 : value = 'h288B;    //value='d10379;             
          'd1655 : value = 'h2891;    //value='d10385;             
          'd1656 : value = 'h2896;    //value='d10390;             
          'd1657 : value = 'h289C;    //value='d10396;             
          'd1658 : value = 'h28A2;    //value='d10402;             
          'd1659 : value = 'h28A8;    //value='d10408;             
          'd1660 : value = 'h28AE;    //value='d10414;             
          'd1661 : value = 'h28B4;    //value='d10420;             
          'd1662 : value = 'h28BA;    //value='d10426;             
          'd1663 : value = 'h28BF;    //value='d10431;             
          'd1664 : value = 'h28C5;    //value='d10437;             
          'd1665 : value = 'h28CB;    //value='d10443;             
          'd1666 : value = 'h28D1;    //value='d10449;             
          'd1667 : value = 'h28D7;    //value='d10455;             
          'd1668 : value = 'h28DD;    //value='d10461;             
          'd1669 : value = 'h28E3;    //value='d10467;             
          'd1670 : value = 'h28E9;    //value='d10473;             
          'd1671 : value = 'h28EE;    //value='d10478;             
          'd1672 : value = 'h28F4;    //value='d10484;             
          'd1673 : value = 'h28FA;    //value='d10490;             
          'd1674 : value = 'h2900;    //value='d10496;             
          'd1675 : value = 'h2906;    //value='d10502;             
          'd1676 : value = 'h290C;    //value='d10508;             
          'd1677 : value = 'h2912;    //value='d10514;             
          'd1678 : value = 'h2918;    //value='d10520;             
          'd1679 : value = 'h291E;    //value='d10526;             
          'd1680 : value = 'h2924;    //value='d10532;             
          'd1681 : value = 'h292A;    //value='d10538;             
          'd1682 : value = 'h292F;    //value='d10543;             
          'd1683 : value = 'h2935;    //value='d10549;             
          'd1684 : value = 'h293B;    //value='d10555;             
          'd1685 : value = 'h2941;    //value='d10561;             
          'd1686 : value = 'h2947;    //value='d10567;             
          'd1687 : value = 'h294D;    //value='d10573;             
          'd1688 : value = 'h2953;    //value='d10579;             
          'd1689 : value = 'h2959;    //value='d10585;             
          'd1690 : value = 'h295F;    //value='d10591;             
          'd1691 : value = 'h2965;    //value='d10597;             
          'd1692 : value = 'h296B;    //value='d10603;             
          'd1693 : value = 'h2971;    //value='d10609;             
          'd1694 : value = 'h2977;    //value='d10615;             
          'd1695 : value = 'h297D;    //value='d10621;             
          'd1696 : value = 'h2983;    //value='d10627;             
          'd1697 : value = 'h2989;    //value='d10633;             
          'd1698 : value = 'h298F;    //value='d10639;             
          'd1699 : value = 'h2995;    //value='d10645;             
          'd1700 : value = 'h299B;    //value='d10651;             
          'd1701 : value = 'h29A1;    //value='d10657;             
          'd1702 : value = 'h29A7;    //value='d10663;             
          'd1703 : value = 'h29AD;    //value='d10669;             
          'd1704 : value = 'h29B3;    //value='d10675;             
          'd1705 : value = 'h29B9;    //value='d10681;             
          'd1706 : value = 'h29BF;    //value='d10687;             
          'd1707 : value = 'h29C5;    //value='d10693;             
          'd1708 : value = 'h29CB;    //value='d10699;             
          'd1709 : value = 'h29D1;    //value='d10705;             
          'd1710 : value = 'h29D7;    //value='d10711;             
          'd1711 : value = 'h29DD;    //value='d10717;             
          'd1712 : value = 'h29E3;    //value='d10723;             
          'd1713 : value = 'h29E9;    //value='d10729;             
          'd1714 : value = 'h29EF;    //value='d10735;             
          'd1715 : value = 'h29F5;    //value='d10741;             
          'd1716 : value = 'h29FB;    //value='d10747;             
          'd1717 : value = 'h2A01;    //value='d10753;             
          'd1718 : value = 'h2A07;    //value='d10759;             
          'd1719 : value = 'h2A0D;    //value='d10765;             
          'd1720 : value = 'h2A13;    //value='d10771;             
          'd1721 : value = 'h2A19;    //value='d10777;             
          'd1722 : value = 'h2A1F;    //value='d10783;             
          'd1723 : value = 'h2A25;    //value='d10789;             
          'd1724 : value = 'h2A2B;    //value='d10795;             
          'd1725 : value = 'h2A31;    //value='d10801;             
          'd1726 : value = 'h2A38;    //value='d10808;             
          'd1727 : value = 'h2A3E;    //value='d10814;             
          'd1728 : value = 'h2A44;    //value='d10820;             
          'd1729 : value = 'h2A4A;    //value='d10826;             
          'd1730 : value = 'h2A50;    //value='d10832;             
          'd1731 : value = 'h2A56;    //value='d10838;             
          'd1732 : value = 'h2A5C;    //value='d10844;             
          'd1733 : value = 'h2A62;    //value='d10850;             
          'd1734 : value = 'h2A68;    //value='d10856;             
          'd1735 : value = 'h2A6E;    //value='d10862;             
          'd1736 : value = 'h2A74;    //value='d10868;             
          'd1737 : value = 'h2A7B;    //value='d10875;             
          'd1738 : value = 'h2A81;    //value='d10881;             
          'd1739 : value = 'h2A87;    //value='d10887;             
          'd1740 : value = 'h2A8D;    //value='d10893;             
          'd1741 : value = 'h2A93;    //value='d10899;             
          'd1742 : value = 'h2A99;    //value='d10905;             
          'd1743 : value = 'h2A9F;    //value='d10911;             
          'd1744 : value = 'h2AA5;    //value='d10917;             
          'd1745 : value = 'h2AAC;    //value='d10924;             
          'd1746 : value = 'h2AB2;    //value='d10930;             
          'd1747 : value = 'h2AB8;    //value='d10936;             
          'd1748 : value = 'h2ABE;    //value='d10942;             
          'd1749 : value = 'h2AC4;    //value='d10948;             
          'd1750 : value = 'h2ACA;    //value='d10954;             
          'd1751 : value = 'h2AD1;    //value='d10961;             
          'd1752 : value = 'h2AD7;    //value='d10967;             
          'd1753 : value = 'h2ADD;    //value='d10973;             
          'd1754 : value = 'h2AE3;    //value='d10979;             
          'd1755 : value = 'h2AE9;    //value='d10985;             
          'd1756 : value = 'h2AEF;    //value='d10991;             
          'd1757 : value = 'h2AF6;    //value='d10998;             
          'd1758 : value = 'h2AFC;    //value='d11004;             
          'd1759 : value = 'h2B02;    //value='d11010;             
          'd1760 : value = 'h2B08;    //value='d11016;             
          'd1761 : value = 'h2B0E;    //value='d11022;             
          'd1762 : value = 'h2B14;    //value='d11028;             
          'd1763 : value = 'h2B1B;    //value='d11035;             
          'd1764 : value = 'h2B21;    //value='d11041;             
          'd1765 : value = 'h2B27;    //value='d11047;             
          'd1766 : value = 'h2B2D;    //value='d11053;             
          'd1767 : value = 'h2B34;    //value='d11060;             
          'd1768 : value = 'h2B3A;    //value='d11066;             
          'd1769 : value = 'h2B40;    //value='d11072;             
          'd1770 : value = 'h2B46;    //value='d11078;             
          'd1771 : value = 'h2B4C;    //value='d11084;             
          'd1772 : value = 'h2B53;    //value='d11091;             
          'd1773 : value = 'h2B59;    //value='d11097;             
          'd1774 : value = 'h2B5F;    //value='d11103;             
          'd1775 : value = 'h2B65;    //value='d11109;             
          'd1776 : value = 'h2B6C;    //value='d11116;             
          'd1777 : value = 'h2B72;    //value='d11122;             
          'd1778 : value = 'h2B78;    //value='d11128;             
          'd1779 : value = 'h2B7E;    //value='d11134;             
          'd1780 : value = 'h2B85;    //value='d11141;             
          'd1781 : value = 'h2B8B;    //value='d11147;             
          'd1782 : value = 'h2B91;    //value='d11153;             
          'd1783 : value = 'h2B97;    //value='d11159;             
          'd1784 : value = 'h2B9E;    //value='d11166;             
          'd1785 : value = 'h2BA4;    //value='d11172;             
          'd1786 : value = 'h2BAA;    //value='d11178;             
          'd1787 : value = 'h2BB1;    //value='d11185;             
          'd1788 : value = 'h2BB7;    //value='d11191;             
          'd1789 : value = 'h2BBD;    //value='d11197;             
          'd1790 : value = 'h2BC3;    //value='d11203;             
          'd1791 : value = 'h2BCA;    //value='d11210;             
          'd1792 : value = 'h2BD0;    //value='d11216;             
          'd1793 : value = 'h2BD6;    //value='d11222;             
          'd1794 : value = 'h2BDD;    //value='d11229;             
          'd1795 : value = 'h2BE3;    //value='d11235;             
          'd1796 : value = 'h2BE9;    //value='d11241;             
          'd1797 : value = 'h2BF0;    //value='d11248;             
          'd1798 : value = 'h2BF6;    //value='d11254;             
          'd1799 : value = 'h2BFC;    //value='d11260;             
          'd1800 : value = 'h2C03;    //value='d11267;             
          'd1801 : value = 'h2C09;    //value='d11273;             
          'd1802 : value = 'h2C0F;    //value='d11279;             
          'd1803 : value = 'h2C16;    //value='d11286;             
          'd1804 : value = 'h2C1C;    //value='d11292;             
          'd1805 : value = 'h2C22;    //value='d11298;             
          'd1806 : value = 'h2C29;    //value='d11305;             
          'd1807 : value = 'h2C2F;    //value='d11311;             
          'd1808 : value = 'h2C35;    //value='d11317;             
          'd1809 : value = 'h2C3C;    //value='d11324;             
          'd1810 : value = 'h2C42;    //value='d11330;             
          'd1811 : value = 'h2C49;    //value='d11337;             
          'd1812 : value = 'h2C4F;    //value='d11343;             
          'd1813 : value = 'h2C55;    //value='d11349;             
          'd1814 : value = 'h2C5C;    //value='d11356;             
          'd1815 : value = 'h2C62;    //value='d11362;             
          'd1816 : value = 'h2C68;    //value='d11368;             
          'd1817 : value = 'h2C6F;    //value='d11375;             
          'd1818 : value = 'h2C75;    //value='d11381;             
          'd1819 : value = 'h2C7C;    //value='d11388;             
          'd1820 : value = 'h2C82;    //value='d11394;             
          'd1821 : value = 'h2C88;    //value='d11400;             
          'd1822 : value = 'h2C8F;    //value='d11407;             
          'd1823 : value = 'h2C95;    //value='d11413;             
          'd1824 : value = 'h2C9C;    //value='d11420;             
          'd1825 : value = 'h2CA2;    //value='d11426;             
          'd1826 : value = 'h2CA9;    //value='d11433;             
          'd1827 : value = 'h2CAF;    //value='d11439;             
          'd1828 : value = 'h2CB5;    //value='d11445;             
          'd1829 : value = 'h2CBC;    //value='d11452;             
          'd1830 : value = 'h2CC2;    //value='d11458;             
          'd1831 : value = 'h2CC9;    //value='d11465;             
          'd1832 : value = 'h2CCF;    //value='d11471;             
          'd1833 : value = 'h2CD6;    //value='d11478;             
          'd1834 : value = 'h2CDC;    //value='d11484;             
          'd1835 : value = 'h2CE3;    //value='d11491;             
          'd1836 : value = 'h2CE9;    //value='d11497;             
          'd1837 : value = 'h2CEF;    //value='d11503;             
          'd1838 : value = 'h2CF6;    //value='d11510;             
          'd1839 : value = 'h2CFC;    //value='d11516;             
          'd1840 : value = 'h2D03;    //value='d11523;             
          'd1841 : value = 'h2D09;    //value='d11529;             
          'd1842 : value = 'h2D10;    //value='d11536;             
          'd1843 : value = 'h2D16;    //value='d11542;             
          'd1844 : value = 'h2D1D;    //value='d11549;             
          'd1845 : value = 'h2D23;    //value='d11555;             
          'd1846 : value = 'h2D2A;    //value='d11562;             
          'd1847 : value = 'h2D30;    //value='d11568;             
          'd1848 : value = 'h2D37;    //value='d11575;             
          'd1849 : value = 'h2D3D;    //value='d11581;             
          'd1850 : value = 'h2D44;    //value='d11588;             
          'd1851 : value = 'h2D4A;    //value='d11594;             
          'd1852 : value = 'h2D51;    //value='d11601;             
          'd1853 : value = 'h2D57;    //value='d11607;             
          'd1854 : value = 'h2D5E;    //value='d11614;             
          'd1855 : value = 'h2D64;    //value='d11620;             
          'd1856 : value = 'h2D6B;    //value='d11627;             
          'd1857 : value = 'h2D72;    //value='d11634;             
          'd1858 : value = 'h2D78;    //value='d11640;             
          'd1859 : value = 'h2D7F;    //value='d11647;             
          'd1860 : value = 'h2D85;    //value='d11653;             
          'd1861 : value = 'h2D8C;    //value='d11660;             
          'd1862 : value = 'h2D92;    //value='d11666;             
          'd1863 : value = 'h2D99;    //value='d11673;             
          'd1864 : value = 'h2D9F;    //value='d11679;             
          'd1865 : value = 'h2DA6;    //value='d11686;             
          'd1866 : value = 'h2DAD;    //value='d11693;             
          'd1867 : value = 'h2DB3;    //value='d11699;             
          'd1868 : value = 'h2DBA;    //value='d11706;             
          'd1869 : value = 'h2DC0;    //value='d11712;             
          'd1870 : value = 'h2DC7;    //value='d11719;             
          'd1871 : value = 'h2DCD;    //value='d11725;             
          'd1872 : value = 'h2DD4;    //value='d11732;             
          'd1873 : value = 'h2DDB;    //value='d11739;             
          'd1874 : value = 'h2DE1;    //value='d11745;             
          'd1875 : value = 'h2DE8;    //value='d11752;             
          'd1876 : value = 'h2DEE;    //value='d11758;             
          'd1877 : value = 'h2DF5;    //value='d11765;             
          'd1878 : value = 'h2DFC;    //value='d11772;             
          'd1879 : value = 'h2E02;    //value='d11778;             
          'd1880 : value = 'h2E09;    //value='d11785;             
          'd1881 : value = 'h2E10;    //value='d11792;             
          'd1882 : value = 'h2E16;    //value='d11798;             
          'd1883 : value = 'h2E1D;    //value='d11805;             
          'd1884 : value = 'h2E23;    //value='d11811;             
          'd1885 : value = 'h2E2A;    //value='d11818;             
          'd1886 : value = 'h2E31;    //value='d11825;             
          'd1887 : value = 'h2E37;    //value='d11831;             
          'd1888 : value = 'h2E3E;    //value='d11838;             
          'd1889 : value = 'h2E45;    //value='d11845;             
          'd1890 : value = 'h2E4B;    //value='d11851;             
          'd1891 : value = 'h2E52;    //value='d11858;             
          'd1892 : value = 'h2E59;    //value='d11865;             
          'd1893 : value = 'h2E5F;    //value='d11871;             
          'd1894 : value = 'h2E66;    //value='d11878;             
          'd1895 : value = 'h2E6D;    //value='d11885;             
          'd1896 : value = 'h2E73;    //value='d11891;             
          'd1897 : value = 'h2E7A;    //value='d11898;             
          'd1898 : value = 'h2E81;    //value='d11905;             
          'd1899 : value = 'h2E87;    //value='d11911;             
          'd1900 : value = 'h2E8E;    //value='d11918;             
          'd1901 : value = 'h2E95;    //value='d11925;             
          'd1902 : value = 'h2E9C;    //value='d11932;             
          'd1903 : value = 'h2EA2;    //value='d11938;             
          'd1904 : value = 'h2EA9;    //value='d11945;             
          'd1905 : value = 'h2EB0;    //value='d11952;             
          'd1906 : value = 'h2EB6;    //value='d11958;             
          'd1907 : value = 'h2EBD;    //value='d11965;             
          'd1908 : value = 'h2EC4;    //value='d11972;             
          'd1909 : value = 'h2ECB;    //value='d11979;             
          'd1910 : value = 'h2ED1;    //value='d11985;             
          'd1911 : value = 'h2ED8;    //value='d11992;             
          'd1912 : value = 'h2EDF;    //value='d11999;             
          'd1913 : value = 'h2EE6;    //value='d12006;             
          'd1914 : value = 'h2EEC;    //value='d12012;             
          'd1915 : value = 'h2EF3;    //value='d12019;             
          'd1916 : value = 'h2EFA;    //value='d12026;             
          'd1917 : value = 'h2F01;    //value='d12033;             
          'd1918 : value = 'h2F07;    //value='d12039;             
          'd1919 : value = 'h2F0E;    //value='d12046;             
          'd1920 : value = 'h2F15;    //value='d12053;             
          'd1921 : value = 'h2F1C;    //value='d12060;             
          'd1922 : value = 'h2F22;    //value='d12066;             
          'd1923 : value = 'h2F29;    //value='d12073;             
          'd1924 : value = 'h2F30;    //value='d12080;             
          'd1925 : value = 'h2F37;    //value='d12087;             
          'd1926 : value = 'h2F3E;    //value='d12094;             
          'd1927 : value = 'h2F44;    //value='d12100;             
          'd1928 : value = 'h2F4B;    //value='d12107;             
          'd1929 : value = 'h2F52;    //value='d12114;             
          'd1930 : value = 'h2F59;    //value='d12121;             
          'd1931 : value = 'h2F60;    //value='d12128;             
          'd1932 : value = 'h2F66;    //value='d12134;             
          'd1933 : value = 'h2F6D;    //value='d12141;             
          'd1934 : value = 'h2F74;    //value='d12148;             
          'd1935 : value = 'h2F7B;    //value='d12155;             
          'd1936 : value = 'h2F82;    //value='d12162;             
          'd1937 : value = 'h2F89;    //value='d12169;             
          'd1938 : value = 'h2F8F;    //value='d12175;             
          'd1939 : value = 'h2F96;    //value='d12182;             
          'd1940 : value = 'h2F9D;    //value='d12189;             
          'd1941 : value = 'h2FA4;    //value='d12196;             
          'd1942 : value = 'h2FAB;    //value='d12203;             
          'd1943 : value = 'h2FB2;    //value='d12210;             
          'd1944 : value = 'h2FB9;    //value='d12217;             
          'd1945 : value = 'h2FC0;    //value='d12224;             
          'd1946 : value = 'h2FC6;    //value='d12230;             
          'd1947 : value = 'h2FCD;    //value='d12237;             
          'd1948 : value = 'h2FD4;    //value='d12244;             
          'd1949 : value = 'h2FDB;    //value='d12251;             
          'd1950 : value = 'h2FE2;    //value='d12258;             
          'd1951 : value = 'h2FE9;    //value='d12265;             
          'd1952 : value = 'h2FF0;    //value='d12272;             
          'd1953 : value = 'h2FF7;    //value='d12279;             
          'd1954 : value = 'h2FFE;    //value='d12286;             
          'd1955 : value = 'h3004;    //value='d12292;             
          'd1956 : value = 'h300B;    //value='d12299;             
          'd1957 : value = 'h3012;    //value='d12306;             
          'd1958 : value = 'h3019;    //value='d12313;             
          'd1959 : value = 'h3020;    //value='d12320;             
          'd1960 : value = 'h3027;    //value='d12327;             
          'd1961 : value = 'h302E;    //value='d12334;             
          'd1962 : value = 'h3035;    //value='d12341;             
          'd1963 : value = 'h303C;    //value='d12348;             
          'd1964 : value = 'h3043;    //value='d12355;             
          'd1965 : value = 'h304A;    //value='d12362;             
          'd1966 : value = 'h3051;    //value='d12369;             
          'd1967 : value = 'h3058;    //value='d12376;             
          'd1968 : value = 'h305F;    //value='d12383;             
          'd1969 : value = 'h3066;    //value='d12390;             
          'd1970 : value = 'h306D;    //value='d12397;             
          'd1971 : value = 'h3073;    //value='d12403;             
          'd1972 : value = 'h307A;    //value='d12410;             
          'd1973 : value = 'h3081;    //value='d12417;             
          'd1974 : value = 'h3088;    //value='d12424;             
          'd1975 : value = 'h308F;    //value='d12431;             
          'd1976 : value = 'h3096;    //value='d12438;             
          'd1977 : value = 'h309D;    //value='d12445;             
          'd1978 : value = 'h30A4;    //value='d12452;             
          'd1979 : value = 'h30AB;    //value='d12459;             
          'd1980 : value = 'h30B2;    //value='d12466;             
          'd1981 : value = 'h30B9;    //value='d12473;             
          'd1982 : value = 'h30C0;    //value='d12480;             
          'd1983 : value = 'h30C7;    //value='d12487;             
          'd1984 : value = 'h30CE;    //value='d12494;             
          'd1985 : value = 'h30D5;    //value='d12501;             
          'd1986 : value = 'h30DD;    //value='d12509;             
          'd1987 : value = 'h30E4;    //value='d12516;             
          'd1988 : value = 'h30EB;    //value='d12523;             
          'd1989 : value = 'h30F2;    //value='d12530;             
          'd1990 : value = 'h30F9;    //value='d12537;             
          'd1991 : value = 'h3100;    //value='d12544;             
          'd1992 : value = 'h3107;    //value='d12551;             
          'd1993 : value = 'h310E;    //value='d12558;             
          'd1994 : value = 'h3115;    //value='d12565;             
          'd1995 : value = 'h311C;    //value='d12572;             
          'd1996 : value = 'h3123;    //value='d12579;             
          'd1997 : value = 'h312A;    //value='d12586;             
          'd1998 : value = 'h3131;    //value='d12593;             
          'd1999 : value = 'h3138;    //value='d12600;             
          'd2000 : value = 'h313F;    //value='d12607;             
          'd2001 : value = 'h3146;    //value='d12614;             
          'd2002 : value = 'h314E;    //value='d12622;             
          'd2003 : value = 'h3155;    //value='d12629;             
          'd2004 : value = 'h315C;    //value='d12636;             
          'd2005 : value = 'h3163;    //value='d12643;             
          'd2006 : value = 'h316A;    //value='d12650;             
          'd2007 : value = 'h3171;    //value='d12657;             
          'd2008 : value = 'h3178;    //value='d12664;             
          'd2009 : value = 'h317F;    //value='d12671;             
          'd2010 : value = 'h3186;    //value='d12678;             
          'd2011 : value = 'h318E;    //value='d12686;             
          'd2012 : value = 'h3195;    //value='d12693;             
          'd2013 : value = 'h319C;    //value='d12700;             
          'd2014 : value = 'h31A3;    //value='d12707;             
          'd2015 : value = 'h31AA;    //value='d12714;             
          'd2016 : value = 'h31B1;    //value='d12721;             
          'd2017 : value = 'h31B8;    //value='d12728;             
          'd2018 : value = 'h31C0;    //value='d12736;             
          'd2019 : value = 'h31C7;    //value='d12743;             
          'd2020 : value = 'h31CE;    //value='d12750;             
          'd2021 : value = 'h31D5;    //value='d12757;             
          'd2022 : value = 'h31DC;    //value='d12764;             
          'd2023 : value = 'h31E3;    //value='d12771;             
          'd2024 : value = 'h31EB;    //value='d12779;             
          'd2025 : value = 'h31F2;    //value='d12786;             
          'd2026 : value = 'h31F9;    //value='d12793;             
          'd2027 : value = 'h3200;    //value='d12800;             
          'd2028 : value = 'h3207;    //value='d12807;             
          'd2029 : value = 'h320F;    //value='d12815;             
          'd2030 : value = 'h3216;    //value='d12822;             
          'd2031 : value = 'h321D;    //value='d12829;             
          'd2032 : value = 'h3224;    //value='d12836;             
          'd2033 : value = 'h322B;    //value='d12843;             
          'd2034 : value = 'h3233;    //value='d12851;             
          'd2035 : value = 'h323A;    //value='d12858;             
          'd2036 : value = 'h3241;    //value='d12865;             
          'd2037 : value = 'h3248;    //value='d12872;             
          'd2038 : value = 'h3250;    //value='d12880;             
          'd2039 : value = 'h3257;    //value='d12887;             
          'd2040 : value = 'h325E;    //value='d12894;             
          'd2041 : value = 'h3265;    //value='d12901;             
          'd2042 : value = 'h326D;    //value='d12909;             
          'd2043 : value = 'h3274;    //value='d12916;             
          'd2044 : value = 'h327B;    //value='d12923;             
          'd2045 : value = 'h3282;    //value='d12930;             
          'd2046 : value = 'h328A;    //value='d12938;             
          'd2047 : value = 'h3291;    //value='d12945;             
          'd2048 : value = 'h3298;    //value='d12952;             
          'd2049 : value = 'h329F;    //value='d12959;             
          'd2050 : value = 'h32A7;    //value='d12967;             
          'd2051 : value = 'h32AE;    //value='d12974;             
          'd2052 : value = 'h32B5;    //value='d12981;             
          'd2053 : value = 'h32BD;    //value='d12989;             
          'd2054 : value = 'h32C4;    //value='d12996;             
          'd2055 : value = 'h32CB;    //value='d13003;             
          'd2056 : value = 'h32D3;    //value='d13011;             
          'd2057 : value = 'h32DA;    //value='d13018;             
          'd2058 : value = 'h32E1;    //value='d13025;             
          'd2059 : value = 'h32E9;    //value='d13033;             
          'd2060 : value = 'h32F0;    //value='d13040;             
          'd2061 : value = 'h32F7;    //value='d13047;             
          'd2062 : value = 'h32FF;    //value='d13055;             
          'd2063 : value = 'h3306;    //value='d13062;             
          'd2064 : value = 'h330D;    //value='d13069;             
          'd2065 : value = 'h3315;    //value='d13077;             
          'd2066 : value = 'h331C;    //value='d13084;             
          'd2067 : value = 'h3323;    //value='d13091;             
          'd2068 : value = 'h332B;    //value='d13099;             
          'd2069 : value = 'h3332;    //value='d13106;             
          'd2070 : value = 'h3339;    //value='d13113;             
          'd2071 : value = 'h3341;    //value='d13121;             
          'd2072 : value = 'h3348;    //value='d13128;             
          'd2073 : value = 'h3350;    //value='d13136;             
          'd2074 : value = 'h3357;    //value='d13143;             
          'd2075 : value = 'h335E;    //value='d13150;             
          'd2076 : value = 'h3366;    //value='d13158;             
          'd2077 : value = 'h336D;    //value='d13165;             
          'd2078 : value = 'h3374;    //value='d13172;             
          'd2079 : value = 'h337C;    //value='d13180;             
          'd2080 : value = 'h3383;    //value='d13187;             
          'd2081 : value = 'h338B;    //value='d13195;             
          'd2082 : value = 'h3392;    //value='d13202;             
          'd2083 : value = 'h339A;    //value='d13210;             
          'd2084 : value = 'h33A1;    //value='d13217;             
          'd2085 : value = 'h33A8;    //value='d13224;             
          'd2086 : value = 'h33B0;    //value='d13232;             
          'd2087 : value = 'h33B7;    //value='d13239;             
          'd2088 : value = 'h33BF;    //value='d13247;             
          'd2089 : value = 'h33C6;    //value='d13254;             
          'd2090 : value = 'h33CE;    //value='d13262;             
          'd2091 : value = 'h33D5;    //value='d13269;             
          'd2092 : value = 'h33DD;    //value='d13277;             
          'd2093 : value = 'h33E4;    //value='d13284;             
          'd2094 : value = 'h33EC;    //value='d13292;             
          'd2095 : value = 'h33F3;    //value='d13299;             
          'd2096 : value = 'h33FA;    //value='d13306;             
          'd2097 : value = 'h3402;    //value='d13314;             
          'd2098 : value = 'h3409;    //value='d13321;             
          'd2099 : value = 'h3411;    //value='d13329;             
          'd2100 : value = 'h3418;    //value='d13336;             
          'd2101 : value = 'h3420;    //value='d13344;             
          'd2102 : value = 'h3427;    //value='d13351;             
          'd2103 : value = 'h342F;    //value='d13359;             
          'd2104 : value = 'h3436;    //value='d13366;             
          'd2105 : value = 'h343E;    //value='d13374;             
          'd2106 : value = 'h3445;    //value='d13381;             
          'd2107 : value = 'h344D;    //value='d13389;             
          'd2108 : value = 'h3455;    //value='d13397;             
          'd2109 : value = 'h345C;    //value='d13404;             
          'd2110 : value = 'h3464;    //value='d13412;             
          'd2111 : value = 'h346B;    //value='d13419;             
          'd2112 : value = 'h3473;    //value='d13427;             
          'd2113 : value = 'h347A;    //value='d13434;             
          'd2114 : value = 'h3482;    //value='d13442;             
          'd2115 : value = 'h3489;    //value='d13449;             
          'd2116 : value = 'h3491;    //value='d13457;             
          'd2117 : value = 'h3498;    //value='d13464;             
          'd2118 : value = 'h34A0;    //value='d13472;             
          'd2119 : value = 'h34A8;    //value='d13480;             
          'd2120 : value = 'h34AF;    //value='d13487;             
          'd2121 : value = 'h34B7;    //value='d13495;             
          'd2122 : value = 'h34BE;    //value='d13502;             
          'd2123 : value = 'h34C6;    //value='d13510;             
          'd2124 : value = 'h34CE;    //value='d13518;             
          'd2125 : value = 'h34D5;    //value='d13525;             
          'd2126 : value = 'h34DD;    //value='d13533;             
          'd2127 : value = 'h34E4;    //value='d13540;             
          'd2128 : value = 'h34EC;    //value='d13548;             
          'd2129 : value = 'h34F4;    //value='d13556;             
          'd2130 : value = 'h34FB;    //value='d13563;             
          'd2131 : value = 'h3503;    //value='d13571;             
          'd2132 : value = 'h350A;    //value='d13578;             
          'd2133 : value = 'h3512;    //value='d13586;             
          'd2134 : value = 'h351A;    //value='d13594;             
          'd2135 : value = 'h3521;    //value='d13601;             
          'd2136 : value = 'h3529;    //value='d13609;             
          'd2137 : value = 'h3531;    //value='d13617;             
          'd2138 : value = 'h3538;    //value='d13624;             
          'd2139 : value = 'h3540;    //value='d13632;             
          'd2140 : value = 'h3548;    //value='d13640;             
          'd2141 : value = 'h354F;    //value='d13647;             
          'd2142 : value = 'h3557;    //value='d13655;             
          'd2143 : value = 'h355F;    //value='d13663;             
          'd2144 : value = 'h3566;    //value='d13670;             
          'd2145 : value = 'h356E;    //value='d13678;             
          'd2146 : value = 'h3576;    //value='d13686;             
          'd2147 : value = 'h357D;    //value='d13693;             
          'd2148 : value = 'h3585;    //value='d13701;             
          'd2149 : value = 'h358D;    //value='d13709;             
          'd2150 : value = 'h3595;    //value='d13717;             
          'd2151 : value = 'h359C;    //value='d13724;             
          'd2152 : value = 'h35A4;    //value='d13732;             
          'd2153 : value = 'h35AC;    //value='d13740;             
          'd2154 : value = 'h35B3;    //value='d13747;             
          'd2155 : value = 'h35BB;    //value='d13755;             
          'd2156 : value = 'h35C3;    //value='d13763;             
          'd2157 : value = 'h35CB;    //value='d13771;             
          'd2158 : value = 'h35D2;    //value='d13778;             
          'd2159 : value = 'h35DA;    //value='d13786;             
          'd2160 : value = 'h35E2;    //value='d13794;             
          'd2161 : value = 'h35EA;    //value='d13802;             
          'd2162 : value = 'h35F1;    //value='d13809;             
          'd2163 : value = 'h35F9;    //value='d13817;             
          'd2164 : value = 'h3601;    //value='d13825;             
          'd2165 : value = 'h3609;    //value='d13833;             
          'd2166 : value = 'h3611;    //value='d13841;             
          'd2167 : value = 'h3618;    //value='d13848;             
          'd2168 : value = 'h3620;    //value='d13856;             
          'd2169 : value = 'h3628;    //value='d13864;             
          'd2170 : value = 'h3630;    //value='d13872;             
          'd2171 : value = 'h3637;    //value='d13879;             
          'd2172 : value = 'h363F;    //value='d13887;             
          'd2173 : value = 'h3647;    //value='d13895;             
          'd2174 : value = 'h364F;    //value='d13903;             
          'd2175 : value = 'h3657;    //value='d13911;             
          'd2176 : value = 'h365F;    //value='d13919;             
          'd2177 : value = 'h3666;    //value='d13926;             
          'd2178 : value = 'h366E;    //value='d13934;             
          'd2179 : value = 'h3676;    //value='d13942;             
          'd2180 : value = 'h367E;    //value='d13950;             
          'd2181 : value = 'h3686;    //value='d13958;             
          'd2182 : value = 'h368E;    //value='d13966;             
          'd2183 : value = 'h3695;    //value='d13973;             
          'd2184 : value = 'h369D;    //value='d13981;             
          'd2185 : value = 'h36A5;    //value='d13989;             
          'd2186 : value = 'h36AD;    //value='d13997;             
          'd2187 : value = 'h36B5;    //value='d14005;             
          'd2188 : value = 'h36BD;    //value='d14013;             
          'd2189 : value = 'h36C5;    //value='d14021;             
          'd2190 : value = 'h36CD;    //value='d14029;             
          'd2191 : value = 'h36D4;    //value='d14036;             
          'd2192 : value = 'h36DC;    //value='d14044;             
          'd2193 : value = 'h36E4;    //value='d14052;             
          'd2194 : value = 'h36EC;    //value='d14060;             
          'd2195 : value = 'h36F4;    //value='d14068;             
          'd2196 : value = 'h36FC;    //value='d14076;             
          'd2197 : value = 'h3704;    //value='d14084;             
          'd2198 : value = 'h370C;    //value='d14092;             
          'd2199 : value = 'h3714;    //value='d14100;             
          'd2200 : value = 'h371C;    //value='d14108;             
          'd2201 : value = 'h3724;    //value='d14116;             
          'd2202 : value = 'h372B;    //value='d14123;             
          'd2203 : value = 'h3733;    //value='d14131;             
          'd2204 : value = 'h373B;    //value='d14139;             
          'd2205 : value = 'h3743;    //value='d14147;             
          'd2206 : value = 'h374B;    //value='d14155;             
          'd2207 : value = 'h3753;    //value='d14163;             
          'd2208 : value = 'h375B;    //value='d14171;             
          'd2209 : value = 'h3763;    //value='d14179;             
          'd2210 : value = 'h376B;    //value='d14187;             
          'd2211 : value = 'h3773;    //value='d14195;             
          'd2212 : value = 'h377B;    //value='d14203;             
          'd2213 : value = 'h3783;    //value='d14211;             
          'd2214 : value = 'h378B;    //value='d14219;             
          'd2215 : value = 'h3793;    //value='d14227;             
          'd2216 : value = 'h379B;    //value='d14235;             
          'd2217 : value = 'h37A3;    //value='d14243;             
          'd2218 : value = 'h37AB;    //value='d14251;             
          'd2219 : value = 'h37B3;    //value='d14259;             
          'd2220 : value = 'h37BB;    //value='d14267;             
          'd2221 : value = 'h37C3;    //value='d14275;             
          'd2222 : value = 'h37CB;    //value='d14283;             
          'd2223 : value = 'h37D3;    //value='d14291;             
          'd2224 : value = 'h37DB;    //value='d14299;             
          'd2225 : value = 'h37E3;    //value='d14307;             
          'd2226 : value = 'h37EB;    //value='d14315;             
          'd2227 : value = 'h37F3;    //value='d14323;             
          'd2228 : value = 'h37FB;    //value='d14331;             
          'd2229 : value = 'h3804;    //value='d14340;             
          'd2230 : value = 'h380C;    //value='d14348;             
          'd2231 : value = 'h3814;    //value='d14356;             
          'd2232 : value = 'h381C;    //value='d14364;             
          'd2233 : value = 'h3824;    //value='d14372;             
          'd2234 : value = 'h382C;    //value='d14380;             
          'd2235 : value = 'h3834;    //value='d14388;             
          'd2236 : value = 'h383C;    //value='d14396;             
          'd2237 : value = 'h3844;    //value='d14404;             
          'd2238 : value = 'h384C;    //value='d14412;             
          'd2239 : value = 'h3854;    //value='d14420;             
          'd2240 : value = 'h385C;    //value='d14428;             
          'd2241 : value = 'h3865;    //value='d14437;             
          'd2242 : value = 'h386D;    //value='d14445;             
          'd2243 : value = 'h3875;    //value='d14453;             
          'd2244 : value = 'h387D;    //value='d14461;             
          'd2245 : value = 'h3885;    //value='d14469;             
          'd2246 : value = 'h388D;    //value='d14477;             
          'd2247 : value = 'h3895;    //value='d14485;             
          'd2248 : value = 'h389D;    //value='d14493;             
          'd2249 : value = 'h38A6;    //value='d14502;             
          'd2250 : value = 'h38AE;    //value='d14510;             
          'd2251 : value = 'h38B6;    //value='d14518;             
          'd2252 : value = 'h38BE;    //value='d14526;             
          'd2253 : value = 'h38C6;    //value='d14534;             
          'd2254 : value = 'h38CE;    //value='d14542;             
          'd2255 : value = 'h38D7;    //value='d14551;             
          'd2256 : value = 'h38DF;    //value='d14559;             
          'd2257 : value = 'h38E7;    //value='d14567;             
          'd2258 : value = 'h38EF;    //value='d14575;             
          'd2259 : value = 'h38F7;    //value='d14583;             
          'd2260 : value = 'h3900;    //value='d14592;             
          'd2261 : value = 'h3908;    //value='d14600;             
          'd2262 : value = 'h3910;    //value='d14608;             
          'd2263 : value = 'h3918;    //value='d14616;             
          'd2264 : value = 'h3920;    //value='d14624;             
          'd2265 : value = 'h3929;    //value='d14633;             
          'd2266 : value = 'h3931;    //value='d14641;             
          'd2267 : value = 'h3939;    //value='d14649;             
          'd2268 : value = 'h3941;    //value='d14657;             
          'd2269 : value = 'h394A;    //value='d14666;             
          'd2270 : value = 'h3952;    //value='d14674;             
          'd2271 : value = 'h395A;    //value='d14682;             
          'd2272 : value = 'h3962;    //value='d14690;             
          'd2273 : value = 'h396B;    //value='d14699;             
          'd2274 : value = 'h3973;    //value='d14707;             
          'd2275 : value = 'h397B;    //value='d14715;             
          'd2276 : value = 'h3983;    //value='d14723;             
          'd2277 : value = 'h398C;    //value='d14732;             
          'd2278 : value = 'h3994;    //value='d14740;             
          'd2279 : value = 'h399C;    //value='d14748;             
          'd2280 : value = 'h39A5;    //value='d14757;             
          'd2281 : value = 'h39AD;    //value='d14765;             
          'd2282 : value = 'h39B5;    //value='d14773;             
          'd2283 : value = 'h39BD;    //value='d14781;             
          'd2284 : value = 'h39C6;    //value='d14790;             
          'd2285 : value = 'h39CE;    //value='d14798;             
          'd2286 : value = 'h39D6;    //value='d14806;             
          'd2287 : value = 'h39DF;    //value='d14815;             
          'd2288 : value = 'h39E7;    //value='d14823;             
          'd2289 : value = 'h39EF;    //value='d14831;             
          'd2290 : value = 'h39F8;    //value='d14840;             
          'd2291 : value = 'h3A00;    //value='d14848;             
          'd2292 : value = 'h3A08;    //value='d14856;             
          'd2293 : value = 'h3A11;    //value='d14865;             
          'd2294 : value = 'h3A19;    //value='d14873;             
          'd2295 : value = 'h3A22;    //value='d14882;             
          'd2296 : value = 'h3A2A;    //value='d14890;             
          'd2297 : value = 'h3A32;    //value='d14898;             
          'd2298 : value = 'h3A3B;    //value='d14907;             
          'd2299 : value = 'h3A43;    //value='d14915;             
          'd2300 : value = 'h3A4B;    //value='d14923;             
          'd2301 : value = 'h3A54;    //value='d14932;             
          'd2302 : value = 'h3A5C;    //value='d14940;             
          'd2303 : value = 'h3A65;    //value='d14949;             
          'd2304 : value = 'h3A6D;    //value='d14957;             
          'd2305 : value = 'h3A75;    //value='d14965;             
          'd2306 : value = 'h3A7E;    //value='d14974;             
          'd2307 : value = 'h3A86;    //value='d14982;             
          'd2308 : value = 'h3A8F;    //value='d14991;             
          'd2309 : value = 'h3A97;    //value='d14999;             
          'd2310 : value = 'h3AA0;    //value='d15008;             
          'd2311 : value = 'h3AA8;    //value='d15016;             
          'd2312 : value = 'h3AB0;    //value='d15024;             
          'd2313 : value = 'h3AB9;    //value='d15033;             
          'd2314 : value = 'h3AC1;    //value='d15041;             
          'd2315 : value = 'h3ACA;    //value='d15050;             
          'd2316 : value = 'h3AD2;    //value='d15058;             
          'd2317 : value = 'h3ADB;    //value='d15067;             
          'd2318 : value = 'h3AE3;    //value='d15075;             
          'd2319 : value = 'h3AEC;    //value='d15084;             
          'd2320 : value = 'h3AF4;    //value='d15092;             
          'd2321 : value = 'h3AFD;    //value='d15101;             
          'd2322 : value = 'h3B05;    //value='d15109;             
          'd2323 : value = 'h3B0E;    //value='d15118;             
          'd2324 : value = 'h3B16;    //value='d15126;             
          'd2325 : value = 'h3B1F;    //value='d15135;             
          'd2326 : value = 'h3B27;    //value='d15143;             
          'd2327 : value = 'h3B30;    //value='d15152;             
          'd2328 : value = 'h3B38;    //value='d15160;             
          'd2329 : value = 'h3B41;    //value='d15169;             
          'd2330 : value = 'h3B49;    //value='d15177;             
          'd2331 : value = 'h3B52;    //value='d15186;             
          'd2332 : value = 'h3B5A;    //value='d15194;             
          'd2333 : value = 'h3B63;    //value='d15203;             
          'd2334 : value = 'h3B6B;    //value='d15211;             
          'd2335 : value = 'h3B74;    //value='d15220;             
          'd2336 : value = 'h3B7D;    //value='d15229;             
          'd2337 : value = 'h3B85;    //value='d15237;             
          'd2338 : value = 'h3B8E;    //value='d15246;             
          'd2339 : value = 'h3B96;    //value='d15254;             
          'd2340 : value = 'h3B9F;    //value='d15263;             
          'd2341 : value = 'h3BA7;    //value='d15271;             
          'd2342 : value = 'h3BB0;    //value='d15280;             
          'd2343 : value = 'h3BB9;    //value='d15289;             
          'd2344 : value = 'h3BC1;    //value='d15297;             
          'd2345 : value = 'h3BCA;    //value='d15306;             
          'd2346 : value = 'h3BD2;    //value='d15314;             
          'd2347 : value = 'h3BDB;    //value='d15323;             
          'd2348 : value = 'h3BE4;    //value='d15332;             
          'd2349 : value = 'h3BEC;    //value='d15340;             
          'd2350 : value = 'h3BF5;    //value='d15349;             
          'd2351 : value = 'h3BFD;    //value='d15357;             
          'd2352 : value = 'h3C06;    //value='d15366;             
          'd2353 : value = 'h3C0F;    //value='d15375;             
          'd2354 : value = 'h3C17;    //value='d15383;             
          'd2355 : value = 'h3C20;    //value='d15392;             
          'd2356 : value = 'h3C29;    //value='d15401;             
          'd2357 : value = 'h3C31;    //value='d15409;             
          'd2358 : value = 'h3C3A;    //value='d15418;             
          'd2359 : value = 'h3C43;    //value='d15427;             
          'd2360 : value = 'h3C4B;    //value='d15435;             
          'd2361 : value = 'h3C54;    //value='d15444;             
          'd2362 : value = 'h3C5D;    //value='d15453;             
          'd2363 : value = 'h3C65;    //value='d15461;             
          'd2364 : value = 'h3C6E;    //value='d15470;             
          'd2365 : value = 'h3C77;    //value='d15479;             
          'd2366 : value = 'h3C80;    //value='d15488;             
          'd2367 : value = 'h3C88;    //value='d15496;             
          'd2368 : value = 'h3C91;    //value='d15505;             
          'd2369 : value = 'h3C9A;    //value='d15514;             
          'd2370 : value = 'h3CA2;    //value='d15522;             
          'd2371 : value = 'h3CAB;    //value='d15531;             
          'd2372 : value = 'h3CB4;    //value='d15540;             
          'd2373 : value = 'h3CBD;    //value='d15549;             
          'd2374 : value = 'h3CC5;    //value='d15557;             
          'd2375 : value = 'h3CCE;    //value='d15566;             
          'd2376 : value = 'h3CD7;    //value='d15575;             
          'd2377 : value = 'h3CE0;    //value='d15584;             
          'd2378 : value = 'h3CE8;    //value='d15592;             
          'd2379 : value = 'h3CF1;    //value='d15601;             
          'd2380 : value = 'h3CFA;    //value='d15610;             
          'd2381 : value = 'h3D03;    //value='d15619;             
          'd2382 : value = 'h3D0B;    //value='d15627;             
          'd2383 : value = 'h3D14;    //value='d15636;             
          'd2384 : value = 'h3D1D;    //value='d15645;             
          'd2385 : value = 'h3D26;    //value='d15654;             
          'd2386 : value = 'h3D2F;    //value='d15663;             
          'd2387 : value = 'h3D37;    //value='d15671;             
          'd2388 : value = 'h3D40;    //value='d15680;             
          'd2389 : value = 'h3D49;    //value='d15689;             
          'd2390 : value = 'h3D52;    //value='d15698;             
          'd2391 : value = 'h3D5B;    //value='d15707;             
          'd2392 : value = 'h3D64;    //value='d15716;             
          'd2393 : value = 'h3D6C;    //value='d15724;             
          'd2394 : value = 'h3D75;    //value='d15733;             
          'd2395 : value = 'h3D7E;    //value='d15742;             
          'd2396 : value = 'h3D87;    //value='d15751;             
          'd2397 : value = 'h3D90;    //value='d15760;             
          'd2398 : value = 'h3D99;    //value='d15769;             
          'd2399 : value = 'h3DA2;    //value='d15778;             
          'd2400 : value = 'h3DAA;    //value='d15786;             
          'd2401 : value = 'h3DB3;    //value='d15795;             
          'd2402 : value = 'h3DBC;    //value='d15804;             
          'd2403 : value = 'h3DC5;    //value='d15813;             
          'd2404 : value = 'h3DCE;    //value='d15822;             
          'd2405 : value = 'h3DD7;    //value='d15831;             
          'd2406 : value = 'h3DE0;    //value='d15840;             
          'd2407 : value = 'h3DE9;    //value='d15849;             
          'd2408 : value = 'h3DF2;    //value='d15858;             
          'd2409 : value = 'h3DFA;    //value='d15866;             
          'd2410 : value = 'h3E03;    //value='d15875;             
          'd2411 : value = 'h3E0C;    //value='d15884;             
          'd2412 : value = 'h3E15;    //value='d15893;             
          'd2413 : value = 'h3E1E;    //value='d15902;             
          'd2414 : value = 'h3E27;    //value='d15911;             
          'd2415 : value = 'h3E30;    //value='d15920;             
          'd2416 : value = 'h3E39;    //value='d15929;             
          'd2417 : value = 'h3E42;    //value='d15938;             
          'd2418 : value = 'h3E4B;    //value='d15947;             
          'd2419 : value = 'h3E54;    //value='d15956;             
          'd2420 : value = 'h3E5D;    //value='d15965;             
          'd2421 : value = 'h3E66;    //value='d15974;             
          'd2422 : value = 'h3E6F;    //value='d15983;             
          'd2423 : value = 'h3E78;    //value='d15992;             
          'd2424 : value = 'h3E81;    //value='d16001;             
          'd2425 : value = 'h3E8A;    //value='d16010;             
          'd2426 : value = 'h3E93;    //value='d16019;             
          'd2427 : value = 'h3E9C;    //value='d16028;             
          'd2428 : value = 'h3EA5;    //value='d16037;             
          'd2429 : value = 'h3EAE;    //value='d16046;             
          'd2430 : value = 'h3EB7;    //value='d16055;             
          'd2431 : value = 'h3EC0;    //value='d16064;             
          'd2432 : value = 'h3EC9;    //value='d16073;             
          'd2433 : value = 'h3ED2;    //value='d16082;             
          'd2434 : value = 'h3EDB;    //value='d16091;             
          'd2435 : value = 'h3EE4;    //value='d16100;             
          'd2436 : value = 'h3EED;    //value='d16109;             
          'd2437 : value = 'h3EF6;    //value='d16118;             
          'd2438 : value = 'h3EFF;    //value='d16127;             
          'd2439 : value = 'h3F08;    //value='d16136;             
          'd2440 : value = 'h3F11;    //value='d16145;             
          'd2441 : value = 'h3F1B;    //value='d16155;             
          'd2442 : value = 'h3F24;    //value='d16164;             
          'd2443 : value = 'h3F2D;    //value='d16173;             
          'd2444 : value = 'h3F36;    //value='d16182;             
          'd2445 : value = 'h3F3F;    //value='d16191;             
          'd2446 : value = 'h3F48;    //value='d16200;             
          'd2447 : value = 'h3F51;    //value='d16209;             
          'd2448 : value = 'h3F5A;    //value='d16218;             
          'd2449 : value = 'h3F63;    //value='d16227;             
          'd2450 : value = 'h3F6C;    //value='d16236;             
          'd2451 : value = 'h3F76;    //value='d16246;             
          'd2452 : value = 'h3F7F;    //value='d16255;             
          'd2453 : value = 'h3F88;    //value='d16264;             
          'd2454 : value = 'h3F91;    //value='d16273;             
          'd2455 : value = 'h3F9A;    //value='d16282;             
          'd2456 : value = 'h3FA3;    //value='d16291;             
          'd2457 : value = 'h3FAC;    //value='d16300;             
          'd2458 : value = 'h3FB6;    //value='d16310;             
          'd2459 : value = 'h3FBF;    //value='d16319;             
          'd2460 : value = 'h3FC8;    //value='d16328;             
          'd2461 : value = 'h3FD1;    //value='d16337;             
          'd2462 : value = 'h3FDA;    //value='d16346;             
          'd2463 : value = 'h3FE4;    //value='d16356;             
          'd2464 : value = 'h3FED;    //value='d16365;             
          'd2465 : value = 'h3FF6;    //value='d16374;             
          'd2466 : value = 'h3FFF;    //value='d16383;             
          'd2467 : value = 'h4008;    //value='d16392;             
          'd2468 : value = 'h4012;    //value='d16402;             
          'd2469 : value = 'h401B;    //value='d16411;             
          'd2470 : value = 'h4024;    //value='d16420;             
          'd2471 : value = 'h402D;    //value='d16429;             
          'd2472 : value = 'h4037;    //value='d16439;             
          'd2473 : value = 'h4040;    //value='d16448;             
          'd2474 : value = 'h4049;    //value='d16457;             
          'd2475 : value = 'h4052;    //value='d16466;             
          'd2476 : value = 'h405C;    //value='d16476;             
          'd2477 : value = 'h4065;    //value='d16485;             
          'd2478 : value = 'h406E;    //value='d16494;             
          'd2479 : value = 'h4077;    //value='d16503;             
          'd2480 : value = 'h4081;    //value='d16513;             
          'd2481 : value = 'h408A;    //value='d16522;             
          'd2482 : value = 'h4093;    //value='d16531;             
          'd2483 : value = 'h409C;    //value='d16540;             
          'd2484 : value = 'h40A6;    //value='d16550;             
          'd2485 : value = 'h40AF;    //value='d16559;             
          'd2486 : value = 'h40B8;    //value='d16568;             
          'd2487 : value = 'h40C2;    //value='d16578;             
          'd2488 : value = 'h40CB;    //value='d16587;             
          'd2489 : value = 'h40D4;    //value='d16596;             
          'd2490 : value = 'h40DE;    //value='d16606;             
          'd2491 : value = 'h40E7;    //value='d16615;             
          'd2492 : value = 'h40F0;    //value='d16624;             
          'd2493 : value = 'h40FA;    //value='d16634;             
          'd2494 : value = 'h4103;    //value='d16643;             
          'd2495 : value = 'h410C;    //value='d16652;             
          'd2496 : value = 'h4116;    //value='d16662;             
          'd2497 : value = 'h411F;    //value='d16671;             
          'd2498 : value = 'h4129;    //value='d16681;             
          'd2499 : value = 'h4132;    //value='d16690;             
          'd2500 : value = 'h413B;    //value='d16699;             
          'd2501 : value = 'h4145;    //value='d16709;             
          'd2502 : value = 'h414E;    //value='d16718;             
          'd2503 : value = 'h4157;    //value='d16727;             
          'd2504 : value = 'h4161;    //value='d16737;             
          'd2505 : value = 'h416A;    //value='d16746;             
          'd2506 : value = 'h4174;    //value='d16756;             
          'd2507 : value = 'h417D;    //value='d16765;             
          'd2508 : value = 'h4187;    //value='d16775;             
          'd2509 : value = 'h4190;    //value='d16784;             
          'd2510 : value = 'h4199;    //value='d16793;             
          'd2511 : value = 'h41A3;    //value='d16803;             
          'd2512 : value = 'h41AC;    //value='d16812;             
          'd2513 : value = 'h41B6;    //value='d16822;             
          'd2514 : value = 'h41BF;    //value='d16831;             
          'd2515 : value = 'h41C9;    //value='d16841;             
          'd2516 : value = 'h41D2;    //value='d16850;             
          'd2517 : value = 'h41DC;    //value='d16860;             
          'd2518 : value = 'h41E5;    //value='d16869;             
          'd2519 : value = 'h41EF;    //value='d16879;             
          'd2520 : value = 'h41F8;    //value='d16888;             
          'd2521 : value = 'h4202;    //value='d16898;             
          'd2522 : value = 'h420B;    //value='d16907;             
          'd2523 : value = 'h4215;    //value='d16917;             
          'd2524 : value = 'h421E;    //value='d16926;             
          'd2525 : value = 'h4228;    //value='d16936;             
          'd2526 : value = 'h4231;    //value='d16945;             
          'd2527 : value = 'h423B;    //value='d16955;             
          'd2528 : value = 'h4244;    //value='d16964;             
          'd2529 : value = 'h424E;    //value='d16974;             
          'd2530 : value = 'h4257;    //value='d16983;             
          'd2531 : value = 'h4261;    //value='d16993;             
          'd2532 : value = 'h426A;    //value='d17002;             
          'd2533 : value = 'h4274;    //value='d17012;             
          'd2534 : value = 'h427E;    //value='d17022;             
          'd2535 : value = 'h4287;    //value='d17031;             
          'd2536 : value = 'h4291;    //value='d17041;             
          'd2537 : value = 'h429A;    //value='d17050;             
          'd2538 : value = 'h42A4;    //value='d17060;             
          'd2539 : value = 'h42AD;    //value='d17069;             
          'd2540 : value = 'h42B7;    //value='d17079;             
          'd2541 : value = 'h42C1;    //value='d17089;             
          'd2542 : value = 'h42CA;    //value='d17098;             
          'd2543 : value = 'h42D4;    //value='d17108;             
          'd2544 : value = 'h42DE;    //value='d17118;             
          'd2545 : value = 'h42E7;    //value='d17127;             
          'd2546 : value = 'h42F1;    //value='d17137;             
          'd2547 : value = 'h42FA;    //value='d17146;             
          'd2548 : value = 'h4304;    //value='d17156;             
          'd2549 : value = 'h430E;    //value='d17166;             
          'd2550 : value = 'h4317;    //value='d17175;             
          'd2551 : value = 'h4321;    //value='d17185;             
          'd2552 : value = 'h432B;    //value='d17195;             
          'd2553 : value = 'h4334;    //value='d17204;             
          'd2554 : value = 'h433E;    //value='d17214;             
          'd2555 : value = 'h4348;    //value='d17224;             
          'd2556 : value = 'h4351;    //value='d17233;             
          'd2557 : value = 'h435B;    //value='d17243;             
          'd2558 : value = 'h4365;    //value='d17253;             
          'd2559 : value = 'h436E;    //value='d17262;             
          'd2560 : value = 'h4378;    //value='d17272;             
          'd2561 : value = 'h4382;    //value='d17282;             
          'd2562 : value = 'h438C;    //value='d17292;             
          'd2563 : value = 'h4395;    //value='d17301;             
          'd2564 : value = 'h439F;    //value='d17311;             
          'd2565 : value = 'h43A9;    //value='d17321;             
          'd2566 : value = 'h43B3;    //value='d17331;             
          'd2567 : value = 'h43BC;    //value='d17340;             
          'd2568 : value = 'h43C6;    //value='d17350;             
          'd2569 : value = 'h43D0;    //value='d17360;             
          'd2570 : value = 'h43DA;    //value='d17370;             
          'd2571 : value = 'h43E3;    //value='d17379;             
          'd2572 : value = 'h43ED;    //value='d17389;             
          'd2573 : value = 'h43F7;    //value='d17399;             
          'd2574 : value = 'h4401;    //value='d17409;             
          'd2575 : value = 'h440A;    //value='d17418;             
          'd2576 : value = 'h4414;    //value='d17428;             
          'd2577 : value = 'h441E;    //value='d17438;             
          'd2578 : value = 'h4428;    //value='d17448;             
          'd2579 : value = 'h4432;    //value='d17458;             
          'd2580 : value = 'h443B;    //value='d17467;             
          'd2581 : value = 'h4445;    //value='d17477;             
          'd2582 : value = 'h444F;    //value='d17487;             
          'd2583 : value = 'h4459;    //value='d17497;             
          'd2584 : value = 'h4463;    //value='d17507;             
          'd2585 : value = 'h446D;    //value='d17517;             
          'd2586 : value = 'h4477;    //value='d17527;             
          'd2587 : value = 'h4480;    //value='d17536;             
          'd2588 : value = 'h448A;    //value='d17546;             
          'd2589 : value = 'h4494;    //value='d17556;             
          'd2590 : value = 'h449E;    //value='d17566;             
          'd2591 : value = 'h44A8;    //value='d17576;             
          'd2592 : value = 'h44B2;    //value='d17586;             
          'd2593 : value = 'h44BC;    //value='d17596;             
          'd2594 : value = 'h44C6;    //value='d17606;             
          'd2595 : value = 'h44CF;    //value='d17615;             
          'd2596 : value = 'h44D9;    //value='d17625;             
          'd2597 : value = 'h44E3;    //value='d17635;             
          'd2598 : value = 'h44ED;    //value='d17645;             
          'd2599 : value = 'h44F7;    //value='d17655;             
          'd2600 : value = 'h4501;    //value='d17665;             
          'd2601 : value = 'h450B;    //value='d17675;             
          'd2602 : value = 'h4515;    //value='d17685;             
          'd2603 : value = 'h451F;    //value='d17695;             
          'd2604 : value = 'h4529;    //value='d17705;             
          'd2605 : value = 'h4533;    //value='d17715;             
          'd2606 : value = 'h453D;    //value='d17725;             
          'd2607 : value = 'h4547;    //value='d17735;             
          'd2608 : value = 'h4551;    //value='d17745;             
          'd2609 : value = 'h455B;    //value='d17755;             
          'd2610 : value = 'h4565;    //value='d17765;             
          'd2611 : value = 'h456F;    //value='d17775;             
          'd2612 : value = 'h4579;    //value='d17785;             
          'd2613 : value = 'h4583;    //value='d17795;             
          'd2614 : value = 'h458D;    //value='d17805;             
          'd2615 : value = 'h4597;    //value='d17815;             
          'd2616 : value = 'h45A1;    //value='d17825;             
          'd2617 : value = 'h45AB;    //value='d17835;             
          'd2618 : value = 'h45B5;    //value='d17845;             
          'd2619 : value = 'h45BF;    //value='d17855;             
          'd2620 : value = 'h45C9;    //value='d17865;             
          'd2621 : value = 'h45D3;    //value='d17875;             
          'd2622 : value = 'h45DD;    //value='d17885;             
          'd2623 : value = 'h45E7;    //value='d17895;             
          'd2624 : value = 'h45F1;    //value='d17905;             
          'd2625 : value = 'h45FB;    //value='d17915;             
          'd2626 : value = 'h4605;    //value='d17925;             
          'd2627 : value = 'h460F;    //value='d17935;             
          'd2628 : value = 'h4619;    //value='d17945;             
          'd2629 : value = 'h4623;    //value='d17955;             
          'd2630 : value = 'h462D;    //value='d17965;             
          'd2631 : value = 'h4638;    //value='d17976;             
          'd2632 : value = 'h4642;    //value='d17986;             
          'd2633 : value = 'h464C;    //value='d17996;             
          'd2634 : value = 'h4656;    //value='d18006;             
          'd2635 : value = 'h4660;    //value='d18016;             
          'd2636 : value = 'h466A;    //value='d18026;             
          'd2637 : value = 'h4674;    //value='d18036;             
          'd2638 : value = 'h467E;    //value='d18046;             
          'd2639 : value = 'h4689;    //value='d18057;             
          'd2640 : value = 'h4693;    //value='d18067;             
          'd2641 : value = 'h469D;    //value='d18077;             
          'd2642 : value = 'h46A7;    //value='d18087;             
          'd2643 : value = 'h46B1;    //value='d18097;             
          'd2644 : value = 'h46BB;    //value='d18107;             
          'd2645 : value = 'h46C6;    //value='d18118;             
          'd2646 : value = 'h46D0;    //value='d18128;             
          'd2647 : value = 'h46DA;    //value='d18138;             
          'd2648 : value = 'h46E4;    //value='d18148;             
          'd2649 : value = 'h46EE;    //value='d18158;             
          'd2650 : value = 'h46F9;    //value='d18169;             
          'd2651 : value = 'h4703;    //value='d18179;             
          'd2652 : value = 'h470D;    //value='d18189;             
          'd2653 : value = 'h4717;    //value='d18199;             
          'd2654 : value = 'h4721;    //value='d18209;             
          'd2655 : value = 'h472C;    //value='d18220;             
          'd2656 : value = 'h4736;    //value='d18230;             
          'd2657 : value = 'h4740;    //value='d18240;             
          'd2658 : value = 'h474A;    //value='d18250;             
          'd2659 : value = 'h4755;    //value='d18261;             
          'd2660 : value = 'h475F;    //value='d18271;             
          'd2661 : value = 'h4769;    //value='d18281;             
          'd2662 : value = 'h4774;    //value='d18292;             
          'd2663 : value = 'h477E;    //value='d18302;             
          'd2664 : value = 'h4788;    //value='d18312;             
          'd2665 : value = 'h4792;    //value='d18322;             
          'd2666 : value = 'h479D;    //value='d18333;             
          'd2667 : value = 'h47A7;    //value='d18343;             
          'd2668 : value = 'h47B1;    //value='d18353;             
          'd2669 : value = 'h47BC;    //value='d18364;             
          'd2670 : value = 'h47C6;    //value='d18374;             
          'd2671 : value = 'h47D0;    //value='d18384;             
          'd2672 : value = 'h47DB;    //value='d18395;             
          'd2673 : value = 'h47E5;    //value='d18405;             
          'd2674 : value = 'h47EF;    //value='d18415;             
          'd2675 : value = 'h47FA;    //value='d18426;             
          'd2676 : value = 'h4804;    //value='d18436;             
          'd2677 : value = 'h480E;    //value='d18446;             
          'd2678 : value = 'h4819;    //value='d18457;             
          'd2679 : value = 'h4823;    //value='d18467;             
          'd2680 : value = 'h482E;    //value='d18478;             
          'd2681 : value = 'h4838;    //value='d18488;             
          'd2682 : value = 'h4842;    //value='d18498;             
          'd2683 : value = 'h484D;    //value='d18509;             
          'd2684 : value = 'h4857;    //value='d18519;             
          'd2685 : value = 'h4862;    //value='d18530;             
          'd2686 : value = 'h486C;    //value='d18540;             
          'd2687 : value = 'h4876;    //value='d18550;             
          'd2688 : value = 'h4881;    //value='d18561;             
          'd2689 : value = 'h488B;    //value='d18571;             
          'd2690 : value = 'h4896;    //value='d18582;             
          'd2691 : value = 'h48A0;    //value='d18592;             
          'd2692 : value = 'h48AB;    //value='d18603;             
          'd2693 : value = 'h48B5;    //value='d18613;             
          'd2694 : value = 'h48C0;    //value='d18624;             
          'd2695 : value = 'h48CA;    //value='d18634;             
          'd2696 : value = 'h48D5;    //value='d18645;             
          'd2697 : value = 'h48DF;    //value='d18655;             
          'd2698 : value = 'h48EA;    //value='d18666;             
          'd2699 : value = 'h48F4;    //value='d18676;             
          'd2700 : value = 'h48FF;    //value='d18687;             
          'd2701 : value = 'h4909;    //value='d18697;             
          'd2702 : value = 'h4914;    //value='d18708;             
          'd2703 : value = 'h491E;    //value='d18718;             
          'd2704 : value = 'h4929;    //value='d18729;             
          'd2705 : value = 'h4933;    //value='d18739;             
          'd2706 : value = 'h493E;    //value='d18750;             
          'd2707 : value = 'h4948;    //value='d18760;             
          'd2708 : value = 'h4953;    //value='d18771;             
          'd2709 : value = 'h495D;    //value='d18781;             
          'd2710 : value = 'h4968;    //value='d18792;             
          'd2711 : value = 'h4972;    //value='d18802;             
          'd2712 : value = 'h497D;    //value='d18813;             
          'd2713 : value = 'h4988;    //value='d18824;             
          'd2714 : value = 'h4992;    //value='d18834;             
          'd2715 : value = 'h499D;    //value='d18845;             
          'd2716 : value = 'h49A7;    //value='d18855;             
          'd2717 : value = 'h49B2;    //value='d18866;             
          'd2718 : value = 'h49BD;    //value='d18877;             
          'd2719 : value = 'h49C7;    //value='d18887;             
          'd2720 : value = 'h49D2;    //value='d18898;             
          'd2721 : value = 'h49DC;    //value='d18908;             
          'd2722 : value = 'h49E7;    //value='d18919;             
          'd2723 : value = 'h49F2;    //value='d18930;             
          'd2724 : value = 'h49FC;    //value='d18940;             
          'd2725 : value = 'h4A07;    //value='d18951;             
          'd2726 : value = 'h4A12;    //value='d18962;             
          'd2727 : value = 'h4A1C;    //value='d18972;             
          'd2728 : value = 'h4A27;    //value='d18983;             
          'd2729 : value = 'h4A32;    //value='d18994;             
          'd2730 : value = 'h4A3C;    //value='d19004;             
          'd2731 : value = 'h4A47;    //value='d19015;             
          'd2732 : value = 'h4A52;    //value='d19026;             
          'd2733 : value = 'h4A5C;    //value='d19036;             
          'd2734 : value = 'h4A67;    //value='d19047;             
          'd2735 : value = 'h4A72;    //value='d19058;             
          'd2736 : value = 'h4A7D;    //value='d19069;             
          'd2737 : value = 'h4A87;    //value='d19079;             
          'd2738 : value = 'h4A92;    //value='d19090;             
          'd2739 : value = 'h4A9D;    //value='d19101;             
          'd2740 : value = 'h4AA7;    //value='d19111;             
          'd2741 : value = 'h4AB2;    //value='d19122;             
          'd2742 : value = 'h4ABD;    //value='d19133;             
          'd2743 : value = 'h4AC8;    //value='d19144;             
          'd2744 : value = 'h4AD2;    //value='d19154;             
          'd2745 : value = 'h4ADD;    //value='d19165;             
          'd2746 : value = 'h4AE8;    //value='d19176;             
          'd2747 : value = 'h4AF3;    //value='d19187;             
          'd2748 : value = 'h4AFE;    //value='d19198;             
          'd2749 : value = 'h4B08;    //value='d19208;             
          'd2750 : value = 'h4B13;    //value='d19219;             
          'd2751 : value = 'h4B1E;    //value='d19230;             
          'd2752 : value = 'h4B29;    //value='d19241;             
          'd2753 : value = 'h4B34;    //value='d19252;             
          'd2754 : value = 'h4B3E;    //value='d19262;             
          'd2755 : value = 'h4B49;    //value='d19273;             
          'd2756 : value = 'h4B54;    //value='d19284;             
          'd2757 : value = 'h4B5F;    //value='d19295;             
          'd2758 : value = 'h4B6A;    //value='d19306;             
          'd2759 : value = 'h4B75;    //value='d19317;             
          'd2760 : value = 'h4B80;    //value='d19328;             
          'd2761 : value = 'h4B8A;    //value='d19338;             
          'd2762 : value = 'h4B95;    //value='d19349;             
          'd2763 : value = 'h4BA0;    //value='d19360;             
          'd2764 : value = 'h4BAB;    //value='d19371;             
          'd2765 : value = 'h4BB6;    //value='d19382;             
          'd2766 : value = 'h4BC1;    //value='d19393;             
          'd2767 : value = 'h4BCC;    //value='d19404;             
          'd2768 : value = 'h4BD7;    //value='d19415;             
          'd2769 : value = 'h4BE2;    //value='d19426;             
          'd2770 : value = 'h4BED;    //value='d19437;             
          'd2771 : value = 'h4BF7;    //value='d19447;             
          'd2772 : value = 'h4C02;    //value='d19458;             
          'd2773 : value = 'h4C0D;    //value='d19469;             
          'd2774 : value = 'h4C18;    //value='d19480;             
          'd2775 : value = 'h4C23;    //value='d19491;             
          'd2776 : value = 'h4C2E;    //value='d19502;             
          'd2777 : value = 'h4C39;    //value='d19513;             
          'd2778 : value = 'h4C44;    //value='d19524;             
          'd2779 : value = 'h4C4F;    //value='d19535;             
          'd2780 : value = 'h4C5A;    //value='d19546;             
          'd2781 : value = 'h4C65;    //value='d19557;             
          'd2782 : value = 'h4C70;    //value='d19568;             
          'd2783 : value = 'h4C7B;    //value='d19579;             
          'd2784 : value = 'h4C86;    //value='d19590;             
          'd2785 : value = 'h4C91;    //value='d19601;             
          'd2786 : value = 'h4C9C;    //value='d19612;             
          'd2787 : value = 'h4CA7;    //value='d19623;             
          'd2788 : value = 'h4CB2;    //value='d19634;             
          'd2789 : value = 'h4CBD;    //value='d19645;             
          'd2790 : value = 'h4CC8;    //value='d19656;             
          'd2791 : value = 'h4CD3;    //value='d19667;             
          'd2792 : value = 'h4CDE;    //value='d19678;             
          'd2793 : value = 'h4CE9;    //value='d19689;             
          'd2794 : value = 'h4CF5;    //value='d19701;             
          'd2795 : value = 'h4D00;    //value='d19712;             
          'd2796 : value = 'h4D0B;    //value='d19723;             
          'd2797 : value = 'h4D16;    //value='d19734;             
          'd2798 : value = 'h4D21;    //value='d19745;             
          'd2799 : value = 'h4D2C;    //value='d19756;             
          'd2800 : value = 'h4D37;    //value='d19767;             
          'd2801 : value = 'h4D42;    //value='d19778;             
          'd2802 : value = 'h4D4D;    //value='d19789;             
          'd2803 : value = 'h4D58;    //value='d19800;             
          'd2804 : value = 'h4D64;    //value='d19812;             
          'd2805 : value = 'h4D6F;    //value='d19823;             
          'd2806 : value = 'h4D7A;    //value='d19834;             
          'd2807 : value = 'h4D85;    //value='d19845;             
          'd2808 : value = 'h4D90;    //value='d19856;             
          'd2809 : value = 'h4D9B;    //value='d19867;             
          'd2810 : value = 'h4DA7;    //value='d19879;             
          'd2811 : value = 'h4DB2;    //value='d19890;             
          'd2812 : value = 'h4DBD;    //value='d19901;             
          'd2813 : value = 'h4DC8;    //value='d19912;             
          'd2814 : value = 'h4DD3;    //value='d19923;             
          'd2815 : value = 'h4DDE;    //value='d19934;             
          'd2816 : value = 'h4DEA;    //value='d19946;             
          'd2817 : value = 'h4DF5;    //value='d19957;             
          'd2818 : value = 'h4E00;    //value='d19968;             
          'd2819 : value = 'h4E0B;    //value='d19979;             
          'd2820 : value = 'h4E17;    //value='d19991;             
          'd2821 : value = 'h4E22;    //value='d20002;             
          'd2822 : value = 'h4E2D;    //value='d20013;             
          'd2823 : value = 'h4E38;    //value='d20024;             
          'd2824 : value = 'h4E44;    //value='d20036;             
          'd2825 : value = 'h4E4F;    //value='d20047;             
          'd2826 : value = 'h4E5A;    //value='d20058;             
          'd2827 : value = 'h4E65;    //value='d20069;             
          'd2828 : value = 'h4E71;    //value='d20081;             
          'd2829 : value = 'h4E7C;    //value='d20092;             
          'd2830 : value = 'h4E87;    //value='d20103;             
          'd2831 : value = 'h4E93;    //value='d20115;             
          'd2832 : value = 'h4E9E;    //value='d20126;             
          'd2833 : value = 'h4EA9;    //value='d20137;             
          'd2834 : value = 'h4EB5;    //value='d20149;             
          'd2835 : value = 'h4EC0;    //value='d20160;             
          'd2836 : value = 'h4ECB;    //value='d20171;             
          'd2837 : value = 'h4ED7;    //value='d20183;             
          'd2838 : value = 'h4EE2;    //value='d20194;             
          'd2839 : value = 'h4EED;    //value='d20205;             
          'd2840 : value = 'h4EF9;    //value='d20217;             
          'd2841 : value = 'h4F04;    //value='d20228;             
          'd2842 : value = 'h4F0F;    //value='d20239;             
          'd2843 : value = 'h4F1B;    //value='d20251;             
          'd2844 : value = 'h4F26;    //value='d20262;             
          'd2845 : value = 'h4F32;    //value='d20274;             
          'd2846 : value = 'h4F3D;    //value='d20285;             
          'd2847 : value = 'h4F48;    //value='d20296;             
          'd2848 : value = 'h4F54;    //value='d20308;             
          'd2849 : value = 'h4F5F;    //value='d20319;             
          'd2850 : value = 'h4F6B;    //value='d20331;             
          'd2851 : value = 'h4F76;    //value='d20342;             
          'd2852 : value = 'h4F81;    //value='d20353;             
          'd2853 : value = 'h4F8D;    //value='d20365;             
          'd2854 : value = 'h4F98;    //value='d20376;             
          'd2855 : value = 'h4FA4;    //value='d20388;             
          'd2856 : value = 'h4FAF;    //value='d20399;             
          'd2857 : value = 'h4FBB;    //value='d20411;             
          'd2858 : value = 'h4FC6;    //value='d20422;             
          'd2859 : value = 'h4FD2;    //value='d20434;             
          'd2860 : value = 'h4FDD;    //value='d20445;             
          'd2861 : value = 'h4FE9;    //value='d20457;             
          'd2862 : value = 'h4FF4;    //value='d20468;             
          'd2863 : value = 'h5000;    //value='d20480;             
          'd2864 : value = 'h500B;    //value='d20491;             
          'd2865 : value = 'h5017;    //value='d20503;             
          'd2866 : value = 'h5022;    //value='d20514;             
          'd2867 : value = 'h502E;    //value='d20526;             
          'd2868 : value = 'h5039;    //value='d20537;             
          'd2869 : value = 'h5045;    //value='d20549;             
          'd2870 : value = 'h5050;    //value='d20560;             
          'd2871 : value = 'h505C;    //value='d20572;             
          'd2872 : value = 'h5068;    //value='d20584;             
          'd2873 : value = 'h5073;    //value='d20595;             
          'd2874 : value = 'h507F;    //value='d20607;             
          'd2875 : value = 'h508A;    //value='d20618;             
          'd2876 : value = 'h5096;    //value='d20630;             
          'd2877 : value = 'h50A2;    //value='d20642;             
          'd2878 : value = 'h50AD;    //value='d20653;             
          'd2879 : value = 'h50B9;    //value='d20665;             
          'd2880 : value = 'h50C4;    //value='d20676;             
          'd2881 : value = 'h50D0;    //value='d20688;             
          'd2882 : value = 'h50DC;    //value='d20700;             
          'd2883 : value = 'h50E7;    //value='d20711;             
          'd2884 : value = 'h50F3;    //value='d20723;             
          'd2885 : value = 'h50FF;    //value='d20735;             
          'd2886 : value = 'h510A;    //value='d20746;             
          'd2887 : value = 'h5116;    //value='d20758;             
          'd2888 : value = 'h5122;    //value='d20770;             
          'd2889 : value = 'h512D;    //value='d20781;             
          'd2890 : value = 'h5139;    //value='d20793;             
          'd2891 : value = 'h5145;    //value='d20805;             
          'd2892 : value = 'h5150;    //value='d20816;             
          'd2893 : value = 'h515C;    //value='d20828;             
          'd2894 : value = 'h5168;    //value='d20840;             
          'd2895 : value = 'h5173;    //value='d20851;             
          'd2896 : value = 'h517F;    //value='d20863;             
          'd2897 : value = 'h518B;    //value='d20875;             
          'd2898 : value = 'h5197;    //value='d20887;             
          'd2899 : value = 'h51A2;    //value='d20898;             
          'd2900 : value = 'h51AE;    //value='d20910;             
          'd2901 : value = 'h51BA;    //value='d20922;             
          'd2902 : value = 'h51C6;    //value='d20934;             
          'd2903 : value = 'h51D1;    //value='d20945;             
          'd2904 : value = 'h51DD;    //value='d20957;             
          'd2905 : value = 'h51E9;    //value='d20969;             
          'd2906 : value = 'h51F5;    //value='d20981;             
          'd2907 : value = 'h5201;    //value='d20993;             
          'd2908 : value = 'h520C;    //value='d21004;             
          'd2909 : value = 'h5218;    //value='d21016;             
          'd2910 : value = 'h5224;    //value='d21028;             
          'd2911 : value = 'h5230;    //value='d21040;             
          'd2912 : value = 'h523C;    //value='d21052;             
          'd2913 : value = 'h5248;    //value='d21064;             
          'd2914 : value = 'h5253;    //value='d21075;             
          'd2915 : value = 'h525F;    //value='d21087;             
          'd2916 : value = 'h526B;    //value='d21099;             
          'd2917 : value = 'h5277;    //value='d21111;             
          'd2918 : value = 'h5283;    //value='d21123;             
          'd2919 : value = 'h528F;    //value='d21135;             
          'd2920 : value = 'h529B;    //value='d21147;             
          'd2921 : value = 'h52A6;    //value='d21158;             
          'd2922 : value = 'h52B2;    //value='d21170;             
          'd2923 : value = 'h52BE;    //value='d21182;             
          'd2924 : value = 'h52CA;    //value='d21194;             
          'd2925 : value = 'h52D6;    //value='d21206;             
          'd2926 : value = 'h52E2;    //value='d21218;             
          'd2927 : value = 'h52EE;    //value='d21230;             
          'd2928 : value = 'h52FA;    //value='d21242;             
          'd2929 : value = 'h5306;    //value='d21254;             
          'd2930 : value = 'h5312;    //value='d21266;             
          'd2931 : value = 'h531E;    //value='d21278;             
          'd2932 : value = 'h532A;    //value='d21290;             
          'd2933 : value = 'h5336;    //value='d21302;             
          'd2934 : value = 'h5342;    //value='d21314;             
          'd2935 : value = 'h534E;    //value='d21326;             
          'd2936 : value = 'h535A;    //value='d21338;             
          'd2937 : value = 'h5366;    //value='d21350;             
          'd2938 : value = 'h5372;    //value='d21362;             
          'd2939 : value = 'h537E;    //value='d21374;             
          'd2940 : value = 'h538A;    //value='d21386;             
          'd2941 : value = 'h5396;    //value='d21398;             
          'd2942 : value = 'h53A2;    //value='d21410;             
          'd2943 : value = 'h53AE;    //value='d21422;             
          'd2944 : value = 'h53BA;    //value='d21434;             
          'd2945 : value = 'h53C6;    //value='d21446;             
          'd2946 : value = 'h53D2;    //value='d21458;             
          'd2947 : value = 'h53DE;    //value='d21470;             
          'd2948 : value = 'h53EA;    //value='d21482;             
          'd2949 : value = 'h53F6;    //value='d21494;             
          'd2950 : value = 'h5402;    //value='d21506;             
          'd2951 : value = 'h540E;    //value='d21518;             
          'd2952 : value = 'h541A;    //value='d21530;             
          'd2953 : value = 'h5427;    //value='d21543;             
          'd2954 : value = 'h5433;    //value='d21555;             
          'd2955 : value = 'h543F;    //value='d21567;             
          'd2956 : value = 'h544B;    //value='d21579;             
          'd2957 : value = 'h5457;    //value='d21591;             
          'd2958 : value = 'h5463;    //value='d21603;             
          'd2959 : value = 'h546F;    //value='d21615;             
          'd2960 : value = 'h547B;    //value='d21627;             
          'd2961 : value = 'h5488;    //value='d21640;             
          'd2962 : value = 'h5494;    //value='d21652;             
          'd2963 : value = 'h54A0;    //value='d21664;             
          'd2964 : value = 'h54AC;    //value='d21676;             
          'd2965 : value = 'h54B8;    //value='d21688;             
          'd2966 : value = 'h54C5;    //value='d21701;             
          'd2967 : value = 'h54D1;    //value='d21713;             
          'd2968 : value = 'h54DD;    //value='d21725;             
          'd2969 : value = 'h54E9;    //value='d21737;             
          'd2970 : value = 'h54F5;    //value='d21749;             
          'd2971 : value = 'h5502;    //value='d21762;             
          'd2972 : value = 'h550E;    //value='d21774;             
          'd2973 : value = 'h551A;    //value='d21786;             
          'd2974 : value = 'h5526;    //value='d21798;             
          'd2975 : value = 'h5533;    //value='d21811;             
          'd2976 : value = 'h553F;    //value='d21823;             
          'd2977 : value = 'h554B;    //value='d21835;             
          'd2978 : value = 'h5557;    //value='d21847;             
          'd2979 : value = 'h5564;    //value='d21860;             
          'd2980 : value = 'h5570;    //value='d21872;             
          'd2981 : value = 'h557C;    //value='d21884;             
          'd2982 : value = 'h5589;    //value='d21897;             
          'd2983 : value = 'h5595;    //value='d21909;             
          'd2984 : value = 'h55A1;    //value='d21921;             
          'd2985 : value = 'h55AE;    //value='d21934;             
          'd2986 : value = 'h55BA;    //value='d21946;             
          'd2987 : value = 'h55C6;    //value='d21958;             
          'd2988 : value = 'h55D3;    //value='d21971;             
          'd2989 : value = 'h55DF;    //value='d21983;             
          'd2990 : value = 'h55EB;    //value='d21995;             
          'd2991 : value = 'h55F8;    //value='d22008;             
          'd2992 : value = 'h5604;    //value='d22020;             
          'd2993 : value = 'h5610;    //value='d22032;             
          'd2994 : value = 'h561D;    //value='d22045;             
          'd2995 : value = 'h5629;    //value='d22057;             
          'd2996 : value = 'h5636;    //value='d22070;             
          'd2997 : value = 'h5642;    //value='d22082;             
          'd2998 : value = 'h564E;    //value='d22094;             
          'd2999 : value = 'h565B;    //value='d22107;             
          'd3000 : value = 'h5667;    //value='d22119;             
          'd3001 : value = 'h5674;    //value='d22132;             
          'd3002 : value = 'h5680;    //value='d22144;             
          'd3003 : value = 'h568D;    //value='d22157;             
          'd3004 : value = 'h5699;    //value='d22169;             
          'd3005 : value = 'h56A6;    //value='d22182;             
          'd3006 : value = 'h56B2;    //value='d22194;             
          'd3007 : value = 'h56BF;    //value='d22207;             
          'd3008 : value = 'h56CB;    //value='d22219;             
          'd3009 : value = 'h56D8;    //value='d22232;             
          'd3010 : value = 'h56E4;    //value='d22244;             
          'd3011 : value = 'h56F1;    //value='d22257;             
          'd3012 : value = 'h56FD;    //value='d22269;             
          'd3013 : value = 'h570A;    //value='d22282;             
          'd3014 : value = 'h5716;    //value='d22294;             
          'd3015 : value = 'h5723;    //value='d22307;             
          'd3016 : value = 'h572F;    //value='d22319;             
          'd3017 : value = 'h573C;    //value='d22332;             
          'd3018 : value = 'h5748;    //value='d22344;             
          'd3019 : value = 'h5755;    //value='d22357;             
          'd3020 : value = 'h5761;    //value='d22369;             
          'd3021 : value = 'h576E;    //value='d22382;             
          'd3022 : value = 'h577B;    //value='d22395;             
          'd3023 : value = 'h5787;    //value='d22407;             
          'd3024 : value = 'h5794;    //value='d22420;             
          'd3025 : value = 'h57A0;    //value='d22432;             
          'd3026 : value = 'h57AD;    //value='d22445;             
          'd3027 : value = 'h57BA;    //value='d22458;             
          'd3028 : value = 'h57C6;    //value='d22470;             
          'd3029 : value = 'h57D3;    //value='d22483;             
          'd3030 : value = 'h57E0;    //value='d22496;             
          'd3031 : value = 'h57EC;    //value='d22508;             
          'd3032 : value = 'h57F9;    //value='d22521;             
          'd3033 : value = 'h5806;    //value='d22534;             
          'd3034 : value = 'h5812;    //value='d22546;             
          'd3035 : value = 'h581F;    //value='d22559;             
          'd3036 : value = 'h582C;    //value='d22572;             
          'd3037 : value = 'h5838;    //value='d22584;             
          'd3038 : value = 'h5845;    //value='d22597;             
          'd3039 : value = 'h5852;    //value='d22610;             
          'd3040 : value = 'h585E;    //value='d22622;             
          'd3041 : value = 'h586B;    //value='d22635;             
          'd3042 : value = 'h5878;    //value='d22648;             
          'd3043 : value = 'h5885;    //value='d22661;             
          'd3044 : value = 'h5891;    //value='d22673;             
          'd3045 : value = 'h589E;    //value='d22686;             
          'd3046 : value = 'h58AB;    //value='d22699;             
          'd3047 : value = 'h58B8;    //value='d22712;             
          'd3048 : value = 'h58C4;    //value='d22724;             
          'd3049 : value = 'h58D1;    //value='d22737;             
          'd3050 : value = 'h58DE;    //value='d22750;             
          'd3051 : value = 'h58EB;    //value='d22763;             
          'd3052 : value = 'h58F7;    //value='d22775;             
          'd3053 : value = 'h5904;    //value='d22788;             
          'd3054 : value = 'h5911;    //value='d22801;             
          'd3055 : value = 'h591E;    //value='d22814;             
          'd3056 : value = 'h592B;    //value='d22827;             
          'd3057 : value = 'h5938;    //value='d22840;             
          'd3058 : value = 'h5944;    //value='d22852;             
          'd3059 : value = 'h5951;    //value='d22865;             
          'd3060 : value = 'h595E;    //value='d22878;             
          'd3061 : value = 'h596B;    //value='d22891;             
          'd3062 : value = 'h5978;    //value='d22904;             
          'd3063 : value = 'h5985;    //value='d22917;             
          'd3064 : value = 'h5992;    //value='d22930;             
          'd3065 : value = 'h599F;    //value='d22943;             
          'd3066 : value = 'h59AB;    //value='d22955;             
          'd3067 : value = 'h59B8;    //value='d22968;             
          'd3068 : value = 'h59C5;    //value='d22981;             
          'd3069 : value = 'h59D2;    //value='d22994;             
          'd3070 : value = 'h59DF;    //value='d23007;             
          'd3071 : value = 'h59EC;    //value='d23020;             
          'd3072 : value = 'h59F9;    //value='d23033;             
          'd3073 : value = 'h5A06;    //value='d23046;             
          'd3074 : value = 'h5A13;    //value='d23059;             
          'd3075 : value = 'h5A20;    //value='d23072;             
          'd3076 : value = 'h5A2D;    //value='d23085;             
          'd3077 : value = 'h5A3A;    //value='d23098;             
          'd3078 : value = 'h5A47;    //value='d23111;             
          'd3079 : value = 'h5A54;    //value='d23124;             
          'd3080 : value = 'h5A61;    //value='d23137;             
          'd3081 : value = 'h5A6E;    //value='d23150;             
          'd3082 : value = 'h5A7B;    //value='d23163;             
          'd3083 : value = 'h5A88;    //value='d23176;             
          'd3084 : value = 'h5A95;    //value='d23189;             
          'd3085 : value = 'h5AA2;    //value='d23202;             
          'd3086 : value = 'h5AAF;    //value='d23215;             
          'd3087 : value = 'h5ABC;    //value='d23228;             
          'd3088 : value = 'h5AC9;    //value='d23241;             
          'd3089 : value = 'h5AD6;    //value='d23254;             
          'd3090 : value = 'h5AE3;    //value='d23267;             
          'd3091 : value = 'h5AF0;    //value='d23280;             
          'd3092 : value = 'h5AFD;    //value='d23293;             
          'd3093 : value = 'h5B0B;    //value='d23307;             
          'd3094 : value = 'h5B18;    //value='d23320;             
          'd3095 : value = 'h5B25;    //value='d23333;             
          'd3096 : value = 'h5B32;    //value='d23346;             
          'd3097 : value = 'h5B3F;    //value='d23359;             
          'd3098 : value = 'h5B4C;    //value='d23372;             
          'd3099 : value = 'h5B59;    //value='d23385;             
          'd3100 : value = 'h5B66;    //value='d23398;             
          'd3101 : value = 'h5B74;    //value='d23412;             
          'd3102 : value = 'h5B81;    //value='d23425;             
          'd3103 : value = 'h5B8E;    //value='d23438;             
          'd3104 : value = 'h5B9B;    //value='d23451;             
          'd3105 : value = 'h5BA8;    //value='d23464;             
          'd3106 : value = 'h5BB5;    //value='d23477;             
          'd3107 : value = 'h5BC3;    //value='d23491;             
          'd3108 : value = 'h5BD0;    //value='d23504;             
          'd3109 : value = 'h5BDD;    //value='d23517;             
          'd3110 : value = 'h5BEA;    //value='d23530;             
          'd3111 : value = 'h5BF8;    //value='d23544;             
          'd3112 : value = 'h5C05;    //value='d23557;             
          'd3113 : value = 'h5C12;    //value='d23570;             
          'd3114 : value = 'h5C1F;    //value='d23583;             
          'd3115 : value = 'h5C2D;    //value='d23597;             
          'd3116 : value = 'h5C3A;    //value='d23610;             
          'd3117 : value = 'h5C47;    //value='d23623;             
          'd3118 : value = 'h5C54;    //value='d23636;             
          'd3119 : value = 'h5C62;    //value='d23650;             
          'd3120 : value = 'h5C6F;    //value='d23663;             
          'd3121 : value = 'h5C7C;    //value='d23676;             
          'd3122 : value = 'h5C8A;    //value='d23690;             
          'd3123 : value = 'h5C97;    //value='d23703;             
          'd3124 : value = 'h5CA4;    //value='d23716;             
          'd3125 : value = 'h5CB2;    //value='d23730;             
          'd3126 : value = 'h5CBF;    //value='d23743;             
          'd3127 : value = 'h5CCC;    //value='d23756;             
          'd3128 : value = 'h5CDA;    //value='d23770;             
          'd3129 : value = 'h5CE7;    //value='d23783;             
          'd3130 : value = 'h5CF4;    //value='d23796;             
          'd3131 : value = 'h5D02;    //value='d23810;             
          'd3132 : value = 'h5D0F;    //value='d23823;             
          'd3133 : value = 'h5D1D;    //value='d23837;             
          'd3134 : value = 'h5D2A;    //value='d23850;             
          'd3135 : value = 'h5D37;    //value='d23863;             
          'd3136 : value = 'h5D45;    //value='d23877;             
          'd3137 : value = 'h5D52;    //value='d23890;             
          'd3138 : value = 'h5D60;    //value='d23904;             
          'd3139 : value = 'h5D6D;    //value='d23917;             
          'd3140 : value = 'h5D7B;    //value='d23931;             
          'd3141 : value = 'h5D88;    //value='d23944;             
          'd3142 : value = 'h5D95;    //value='d23957;             
          'd3143 : value = 'h5DA3;    //value='d23971;             
          'd3144 : value = 'h5DB0;    //value='d23984;             
          'd3145 : value = 'h5DBE;    //value='d23998;             
          'd3146 : value = 'h5DCB;    //value='d24011;             
          'd3147 : value = 'h5DD9;    //value='d24025;             
          'd3148 : value = 'h5DE6;    //value='d24038;             
          'd3149 : value = 'h5DF4;    //value='d24052;             
          'd3150 : value = 'h5E01;    //value='d24065;             
          'd3151 : value = 'h5E0F;    //value='d24079;             
          'd3152 : value = 'h5E1D;    //value='d24093;             
          'd3153 : value = 'h5E2A;    //value='d24106;             
          'd3154 : value = 'h5E38;    //value='d24120;             
          'd3155 : value = 'h5E45;    //value='d24133;             
          'd3156 : value = 'h5E53;    //value='d24147;             
          'd3157 : value = 'h5E60;    //value='d24160;             
          'd3158 : value = 'h5E6E;    //value='d24174;             
          'd3159 : value = 'h5E7C;    //value='d24188;             
          'd3160 : value = 'h5E89;    //value='d24201;             
          'd3161 : value = 'h5E97;    //value='d24215;             
          'd3162 : value = 'h5EA4;    //value='d24228;             
          'd3163 : value = 'h5EB2;    //value='d24242;             
          'd3164 : value = 'h5EC0;    //value='d24256;             
          'd3165 : value = 'h5ECD;    //value='d24269;             
          'd3166 : value = 'h5EDB;    //value='d24283;             
          'd3167 : value = 'h5EE9;    //value='d24297;             
          'd3168 : value = 'h5EF6;    //value='d24310;             
          'd3169 : value = 'h5F04;    //value='d24324;             
          'd3170 : value = 'h5F12;    //value='d24338;             
          'd3171 : value = 'h5F1F;    //value='d24351;             
          'd3172 : value = 'h5F2D;    //value='d24365;             
          'd3173 : value = 'h5F3B;    //value='d24379;             
          'd3174 : value = 'h5F48;    //value='d24392;             
          'd3175 : value = 'h5F56;    //value='d24406;             
          'd3176 : value = 'h5F64;    //value='d24420;             
          'd3177 : value = 'h5F72;    //value='d24434;             
          'd3178 : value = 'h5F7F;    //value='d24447;             
          'd3179 : value = 'h5F8D;    //value='d24461;             
          'd3180 : value = 'h5F9B;    //value='d24475;             
          'd3181 : value = 'h5FA9;    //value='d24489;             
          'd3182 : value = 'h5FB6;    //value='d24502;             
          'd3183 : value = 'h5FC4;    //value='d24516;             
          'd3184 : value = 'h5FD2;    //value='d24530;             
          'd3185 : value = 'h5FE0;    //value='d24544;             
          'd3186 : value = 'h5FED;    //value='d24557;             
          'd3187 : value = 'h5FFB;    //value='d24571;             
          'd3188 : value = 'h6009;    //value='d24585;             
          'd3189 : value = 'h6017;    //value='d24599;             
          'd3190 : value = 'h6025;    //value='d24613;             
          'd3191 : value = 'h6033;    //value='d24627;             
          'd3192 : value = 'h6040;    //value='d24640;             
          'd3193 : value = 'h604E;    //value='d24654;             
          'd3194 : value = 'h605C;    //value='d24668;             
          'd3195 : value = 'h606A;    //value='d24682;             
          'd3196 : value = 'h6078;    //value='d24696;             
          'd3197 : value = 'h6086;    //value='d24710;             
          'd3198 : value = 'h6094;    //value='d24724;             
          'd3199 : value = 'h60A2;    //value='d24738;             
          'd3200 : value = 'h60AF;    //value='d24751;             
          'd3201 : value = 'h60BD;    //value='d24765;             
          'd3202 : value = 'h60CB;    //value='d24779;             
          'd3203 : value = 'h60D9;    //value='d24793;             
          'd3204 : value = 'h60E7;    //value='d24807;             
          'd3205 : value = 'h60F5;    //value='d24821;             
          'd3206 : value = 'h6103;    //value='d24835;             
          'd3207 : value = 'h6111;    //value='d24849;             
          'd3208 : value = 'h611F;    //value='d24863;             
          'd3209 : value = 'h612D;    //value='d24877;             
          'd3210 : value = 'h613B;    //value='d24891;             
          'd3211 : value = 'h6149;    //value='d24905;             
          'd3212 : value = 'h6157;    //value='d24919;             
          'd3213 : value = 'h6165;    //value='d24933;             
          'd3214 : value = 'h6173;    //value='d24947;             
          'd3215 : value = 'h6181;    //value='d24961;             
          'd3216 : value = 'h618F;    //value='d24975;             
          'd3217 : value = 'h619D;    //value='d24989;             
          'd3218 : value = 'h61AB;    //value='d25003;             
          'd3219 : value = 'h61B9;    //value='d25017;             
          'd3220 : value = 'h61C7;    //value='d25031;             
          'd3221 : value = 'h61D5;    //value='d25045;             
          'd3222 : value = 'h61E3;    //value='d25059;             
          'd3223 : value = 'h61F2;    //value='d25074;             
          'd3224 : value = 'h6200;    //value='d25088;             
          'd3225 : value = 'h620E;    //value='d25102;             
          'd3226 : value = 'h621C;    //value='d25116;             
          'd3227 : value = 'h622A;    //value='d25130;             
          'd3228 : value = 'h6238;    //value='d25144;             
          'd3229 : value = 'h6246;    //value='d25158;             
          'd3230 : value = 'h6254;    //value='d25172;             
          'd3231 : value = 'h6263;    //value='d25187;             
          'd3232 : value = 'h6271;    //value='d25201;             
          'd3233 : value = 'h627F;    //value='d25215;             
          'd3234 : value = 'h628D;    //value='d25229;             
          'd3235 : value = 'h629B;    //value='d25243;             
          'd3236 : value = 'h62AA;    //value='d25258;             
          'd3237 : value = 'h62B8;    //value='d25272;             
          'd3238 : value = 'h62C6;    //value='d25286;             
          'd3239 : value = 'h62D4;    //value='d25300;             
          'd3240 : value = 'h62E2;    //value='d25314;             
          'd3241 : value = 'h62F1;    //value='d25329;             
          'd3242 : value = 'h62FF;    //value='d25343;             
          'd3243 : value = 'h630D;    //value='d25357;             
          'd3244 : value = 'h631B;    //value='d25371;             
          'd3245 : value = 'h632A;    //value='d25386;             
          'd3246 : value = 'h6338;    //value='d25400;             
          'd3247 : value = 'h6346;    //value='d25414;             
          'd3248 : value = 'h6354;    //value='d25428;             
          'd3249 : value = 'h6363;    //value='d25443;             
          'd3250 : value = 'h6371;    //value='d25457;             
          'd3251 : value = 'h637F;    //value='d25471;             
          'd3252 : value = 'h638E;    //value='d25486;             
          'd3253 : value = 'h639C;    //value='d25500;             
          'd3254 : value = 'h63AA;    //value='d25514;             
          'd3255 : value = 'h63B9;    //value='d25529;             
          'd3256 : value = 'h63C7;    //value='d25543;             
          'd3257 : value = 'h63D5;    //value='d25557;             
          'd3258 : value = 'h63E4;    //value='d25572;             
          'd3259 : value = 'h63F2;    //value='d25586;             
          'd3260 : value = 'h6401;    //value='d25601;             
          'd3261 : value = 'h640F;    //value='d25615;             
          'd3262 : value = 'h641D;    //value='d25629;             
          'd3263 : value = 'h642C;    //value='d25644;             
          'd3264 : value = 'h643A;    //value='d25658;             
          'd3265 : value = 'h6449;    //value='d25673;             
          'd3266 : value = 'h6457;    //value='d25687;             
          'd3267 : value = 'h6466;    //value='d25702;             
          'd3268 : value = 'h6474;    //value='d25716;             
          'd3269 : value = 'h6482;    //value='d25730;             
          'd3270 : value = 'h6491;    //value='d25745;             
          'd3271 : value = 'h649F;    //value='d25759;             
          'd3272 : value = 'h64AE;    //value='d25774;             
          'd3273 : value = 'h64BC;    //value='d25788;             
          'd3274 : value = 'h64CB;    //value='d25803;             
          'd3275 : value = 'h64D9;    //value='d25817;             
          'd3276 : value = 'h64E8;    //value='d25832;             
          'd3277 : value = 'h64F6;    //value='d25846;             
          'd3278 : value = 'h6505;    //value='d25861;             
          'd3279 : value = 'h6513;    //value='d25875;             
          'd3280 : value = 'h6522;    //value='d25890;             
          'd3281 : value = 'h6531;    //value='d25905;             
          'd3282 : value = 'h653F;    //value='d25919;             
          'd3283 : value = 'h654E;    //value='d25934;             
          'd3284 : value = 'h655C;    //value='d25948;             
          'd3285 : value = 'h656B;    //value='d25963;             
          'd3286 : value = 'h657A;    //value='d25978;             
          'd3287 : value = 'h6588;    //value='d25992;             
          'd3288 : value = 'h6597;    //value='d26007;             
          'd3289 : value = 'h65A5;    //value='d26021;             
          'd3290 : value = 'h65B4;    //value='d26036;             
          'd3291 : value = 'h65C3;    //value='d26051;             
          'd3292 : value = 'h65D1;    //value='d26065;             
          'd3293 : value = 'h65E0;    //value='d26080;             
          'd3294 : value = 'h65EF;    //value='d26095;             
          'd3295 : value = 'h65FD;    //value='d26109;             
          'd3296 : value = 'h660C;    //value='d26124;             
          'd3297 : value = 'h661B;    //value='d26139;             
          'd3298 : value = 'h6629;    //value='d26153;             
          'd3299 : value = 'h6638;    //value='d26168;             
          'd3300 : value = 'h6647;    //value='d26183;             
          'd3301 : value = 'h6656;    //value='d26198;             
          'd3302 : value = 'h6664;    //value='d26212;             
          'd3303 : value = 'h6673;    //value='d26227;             
          'd3304 : value = 'h6682;    //value='d26242;             
          'd3305 : value = 'h6690;    //value='d26256;             
          'd3306 : value = 'h669F;    //value='d26271;             
          'd3307 : value = 'h66AE;    //value='d26286;             
          'd3308 : value = 'h66BD;    //value='d26301;             
          'd3309 : value = 'h66CC;    //value='d26316;             
          'd3310 : value = 'h66DA;    //value='d26330;             
          'd3311 : value = 'h66E9;    //value='d26345;             
          'd3312 : value = 'h66F8;    //value='d26360;             
          'd3313 : value = 'h6707;    //value='d26375;             
          'd3314 : value = 'h6716;    //value='d26390;             
          'd3315 : value = 'h6724;    //value='d26404;             
          'd3316 : value = 'h6733;    //value='d26419;             
          'd3317 : value = 'h6742;    //value='d26434;             
          'd3318 : value = 'h6751;    //value='d26449;             
          'd3319 : value = 'h6760;    //value='d26464;             
          'd3320 : value = 'h676F;    //value='d26479;             
          'd3321 : value = 'h677E;    //value='d26494;             
          'd3322 : value = 'h678D;    //value='d26509;             
          'd3323 : value = 'h679C;    //value='d26524;             
          'd3324 : value = 'h67AA;    //value='d26538;             
          'd3325 : value = 'h67B9;    //value='d26553;             
          'd3326 : value = 'h67C8;    //value='d26568;             
          'd3327 : value = 'h67D7;    //value='d26583;             
          'd3328 : value = 'h67E6;    //value='d26598;             
          'd3329 : value = 'h67F5;    //value='d26613;             
          'd3330 : value = 'h6804;    //value='d26628;             
          'd3331 : value = 'h6813;    //value='d26643;             
          'd3332 : value = 'h6822;    //value='d26658;             
          'd3333 : value = 'h6831;    //value='d26673;             
          'd3334 : value = 'h6840;    //value='d26688;             
          'd3335 : value = 'h684F;    //value='d26703;             
          'd3336 : value = 'h685E;    //value='d26718;             
          'd3337 : value = 'h686D;    //value='d26733;             
          'd3338 : value = 'h687C;    //value='d26748;             
          'd3339 : value = 'h688B;    //value='d26763;             
          'd3340 : value = 'h689A;    //value='d26778;             
          'd3341 : value = 'h68A9;    //value='d26793;             
          'd3342 : value = 'h68B8;    //value='d26808;             
          'd3343 : value = 'h68C7;    //value='d26823;             
          'd3344 : value = 'h68D6;    //value='d26838;             
          'd3345 : value = 'h68E6;    //value='d26854;             
          'd3346 : value = 'h68F5;    //value='d26869;             
          'd3347 : value = 'h6904;    //value='d26884;             
          'd3348 : value = 'h6913;    //value='d26899;             
          'd3349 : value = 'h6922;    //value='d26914;             
          'd3350 : value = 'h6931;    //value='d26929;             
          'd3351 : value = 'h6940;    //value='d26944;             
          'd3352 : value = 'h694F;    //value='d26959;             
          'd3353 : value = 'h695F;    //value='d26975;             
          'd3354 : value = 'h696E;    //value='d26990;             
          'd3355 : value = 'h697D;    //value='d27005;             
          'd3356 : value = 'h698C;    //value='d27020;             
          'd3357 : value = 'h699B;    //value='d27035;             
          'd3358 : value = 'h69AB;    //value='d27051;             
          'd3359 : value = 'h69BA;    //value='d27066;             
          'd3360 : value = 'h69C9;    //value='d27081;             
          'd3361 : value = 'h69D8;    //value='d27096;             
          'd3362 : value = 'h69E7;    //value='d27111;             
          'd3363 : value = 'h69F7;    //value='d27127;             
          'd3364 : value = 'h6A06;    //value='d27142;             
          'd3365 : value = 'h6A15;    //value='d27157;             
          'd3366 : value = 'h6A24;    //value='d27172;             
          'd3367 : value = 'h6A34;    //value='d27188;             
          'd3368 : value = 'h6A43;    //value='d27203;             
          'd3369 : value = 'h6A52;    //value='d27218;             
          'd3370 : value = 'h6A62;    //value='d27234;             
          'd3371 : value = 'h6A71;    //value='d27249;             
          'd3372 : value = 'h6A80;    //value='d27264;             
          'd3373 : value = 'h6A90;    //value='d27280;             
          'd3374 : value = 'h6A9F;    //value='d27295;             
          'd3375 : value = 'h6AAE;    //value='d27310;             
          'd3376 : value = 'h6ABE;    //value='d27326;             
          'd3377 : value = 'h6ACD;    //value='d27341;             
          'd3378 : value = 'h6ADC;    //value='d27356;             
          'd3379 : value = 'h6AEC;    //value='d27372;             
          'd3380 : value = 'h6AFB;    //value='d27387;             
          'd3381 : value = 'h6B0B;    //value='d27403;             
          'd3382 : value = 'h6B1A;    //value='d27418;             
          'd3383 : value = 'h6B29;    //value='d27433;             
          'd3384 : value = 'h6B39;    //value='d27449;             
          'd3385 : value = 'h6B48;    //value='d27464;             
          'd3386 : value = 'h6B58;    //value='d27480;             
          'd3387 : value = 'h6B67;    //value='d27495;             
          'd3388 : value = 'h6B77;    //value='d27511;             
          'd3389 : value = 'h6B86;    //value='d27526;             
          'd3390 : value = 'h6B96;    //value='d27542;             
          'd3391 : value = 'h6BA5;    //value='d27557;             
          'd3392 : value = 'h6BB5;    //value='d27573;             
          'd3393 : value = 'h6BC4;    //value='d27588;             
          'd3394 : value = 'h6BD4;    //value='d27604;             
          'd3395 : value = 'h6BE3;    //value='d27619;             
          'd3396 : value = 'h6BF3;    //value='d27635;             
          'd3397 : value = 'h6C02;    //value='d27650;             
          'd3398 : value = 'h6C12;    //value='d27666;             
          'd3399 : value = 'h6C21;    //value='d27681;             
          'd3400 : value = 'h6C31;    //value='d27697;             
          'd3401 : value = 'h6C40;    //value='d27712;             
          'd3402 : value = 'h6C50;    //value='d27728;             
          'd3403 : value = 'h6C60;    //value='d27744;             
          'd3404 : value = 'h6C6F;    //value='d27759;             
          'd3405 : value = 'h6C7F;    //value='d27775;             
          'd3406 : value = 'h6C8E;    //value='d27790;             
          'd3407 : value = 'h6C9E;    //value='d27806;             
          'd3408 : value = 'h6CAE;    //value='d27822;             
          'd3409 : value = 'h6CBD;    //value='d27837;             
          'd3410 : value = 'h6CCD;    //value='d27853;             
          'd3411 : value = 'h6CDD;    //value='d27869;             
          'd3412 : value = 'h6CEC;    //value='d27884;             
          'd3413 : value = 'h6CFC;    //value='d27900;             
          'd3414 : value = 'h6D0C;    //value='d27916;             
          'd3415 : value = 'h6D1B;    //value='d27931;             
          'd3416 : value = 'h6D2B;    //value='d27947;             
          'd3417 : value = 'h6D3B;    //value='d27963;             
          'd3418 : value = 'h6D4B;    //value='d27979;             
          'd3419 : value = 'h6D5A;    //value='d27994;             
          'd3420 : value = 'h6D6A;    //value='d28010;             
          'd3421 : value = 'h6D7A;    //value='d28026;             
          'd3422 : value = 'h6D8A;    //value='d28042;             
          'd3423 : value = 'h6D99;    //value='d28057;             
          'd3424 : value = 'h6DA9;    //value='d28073;             
          'd3425 : value = 'h6DB9;    //value='d28089;             
          'd3426 : value = 'h6DC9;    //value='d28105;             
          'd3427 : value = 'h6DD8;    //value='d28120;             
          'd3428 : value = 'h6DE8;    //value='d28136;             
          'd3429 : value = 'h6DF8;    //value='d28152;             
          'd3430 : value = 'h6E08;    //value='d28168;             
          'd3431 : value = 'h6E18;    //value='d28184;             
          'd3432 : value = 'h6E28;    //value='d28200;             
          'd3433 : value = 'h6E37;    //value='d28215;             
          'd3434 : value = 'h6E47;    //value='d28231;             
          'd3435 : value = 'h6E57;    //value='d28247;             
          'd3436 : value = 'h6E67;    //value='d28263;             
          'd3437 : value = 'h6E77;    //value='d28279;             
          'd3438 : value = 'h6E87;    //value='d28295;             
          'd3439 : value = 'h6E97;    //value='d28311;             
          'd3440 : value = 'h6EA7;    //value='d28327;             
          'd3441 : value = 'h6EB7;    //value='d28343;             
          'd3442 : value = 'h6EC7;    //value='d28359;             
          'd3443 : value = 'h6ED7;    //value='d28375;             
          'd3444 : value = 'h6EE6;    //value='d28390;             
          'd3445 : value = 'h6EF6;    //value='d28406;             
          'd3446 : value = 'h6F06;    //value='d28422;             
          'd3447 : value = 'h6F16;    //value='d28438;             
          'd3448 : value = 'h6F26;    //value='d28454;             
          'd3449 : value = 'h6F36;    //value='d28470;             
          'd3450 : value = 'h6F46;    //value='d28486;             
          'd3451 : value = 'h6F56;    //value='d28502;             
          'd3452 : value = 'h6F66;    //value='d28518;             
          'd3453 : value = 'h6F76;    //value='d28534;             
          'd3454 : value = 'h6F87;    //value='d28551;             
          'd3455 : value = 'h6F97;    //value='d28567;             
          'd3456 : value = 'h6FA7;    //value='d28583;             
          'd3457 : value = 'h6FB7;    //value='d28599;             
          'd3458 : value = 'h6FC7;    //value='d28615;             
          'd3459 : value = 'h6FD7;    //value='d28631;             
          'd3460 : value = 'h6FE7;    //value='d28647;             
          'd3461 : value = 'h6FF7;    //value='d28663;             
          'd3462 : value = 'h7007;    //value='d28679;             
          'd3463 : value = 'h7017;    //value='d28695;             
          'd3464 : value = 'h7027;    //value='d28711;             
          'd3465 : value = 'h7038;    //value='d28728;             
          'd3466 : value = 'h7048;    //value='d28744;             
          'd3467 : value = 'h7058;    //value='d28760;             
          'd3468 : value = 'h7068;    //value='d28776;             
          'd3469 : value = 'h7078;    //value='d28792;             
          'd3470 : value = 'h7088;    //value='d28808;             
          'd3471 : value = 'h7099;    //value='d28825;             
          'd3472 : value = 'h70A9;    //value='d28841;             
          'd3473 : value = 'h70B9;    //value='d28857;             
          'd3474 : value = 'h70C9;    //value='d28873;             
          'd3475 : value = 'h70DA;    //value='d28890;             
          'd3476 : value = 'h70EA;    //value='d28906;             
          'd3477 : value = 'h70FA;    //value='d28922;             
          'd3478 : value = 'h710A;    //value='d28938;             
          'd3479 : value = 'h711B;    //value='d28955;             
          'd3480 : value = 'h712B;    //value='d28971;             
          'd3481 : value = 'h713B;    //value='d28987;             
          'd3482 : value = 'h714B;    //value='d29003;             
          'd3483 : value = 'h715C;    //value='d29020;             
          'd3484 : value = 'h716C;    //value='d29036;             
          'd3485 : value = 'h717C;    //value='d29052;             
          'd3486 : value = 'h718D;    //value='d29069;             
          'd3487 : value = 'h719D;    //value='d29085;             
          'd3488 : value = 'h71AD;    //value='d29101;             
          'd3489 : value = 'h71BE;    //value='d29118;             
          'd3490 : value = 'h71CE;    //value='d29134;             
          'd3491 : value = 'h71DF;    //value='d29151;             
          'd3492 : value = 'h71EF;    //value='d29167;             
          'd3493 : value = 'h71FF;    //value='d29183;             
          'd3494 : value = 'h7210;    //value='d29200;             
          'd3495 : value = 'h7220;    //value='d29216;             
          'd3496 : value = 'h7231;    //value='d29233;             
          'd3497 : value = 'h7241;    //value='d29249;             
          'd3498 : value = 'h7252;    //value='d29266;             
          'd3499 : value = 'h7262;    //value='d29282;             
          'd3500 : value = 'h7272;    //value='d29298;             
          'd3501 : value = 'h7283;    //value='d29315;             
          'd3502 : value = 'h7293;    //value='d29331;             
          'd3503 : value = 'h72A4;    //value='d29348;             
          'd3504 : value = 'h72B4;    //value='d29364;             
          'd3505 : value = 'h72C5;    //value='d29381;             
          'd3506 : value = 'h72D5;    //value='d29397;             
          'd3507 : value = 'h72E6;    //value='d29414;             
          'd3508 : value = 'h72F7;    //value='d29431;             
          'd3509 : value = 'h7307;    //value='d29447;             
          'd3510 : value = 'h7318;    //value='d29464;             
          'd3511 : value = 'h7328;    //value='d29480;             
          'd3512 : value = 'h7339;    //value='d29497;             
          'd3513 : value = 'h7349;    //value='d29513;             
          'd3514 : value = 'h735A;    //value='d29530;             
          'd3515 : value = 'h736B;    //value='d29547;             
          'd3516 : value = 'h737B;    //value='d29563;             
          'd3517 : value = 'h738C;    //value='d29580;             
          'd3518 : value = 'h739C;    //value='d29596;             
          'd3519 : value = 'h73AD;    //value='d29613;             
          'd3520 : value = 'h73BE;    //value='d29630;             
          'd3521 : value = 'h73CE;    //value='d29646;             
          'd3522 : value = 'h73DF;    //value='d29663;             
          'd3523 : value = 'h73F0;    //value='d29680;             
          'd3524 : value = 'h7400;    //value='d29696;             
          'd3525 : value = 'h7411;    //value='d29713;             
          'd3526 : value = 'h7422;    //value='d29730;             
          'd3527 : value = 'h7433;    //value='d29747;             
          'd3528 : value = 'h7443;    //value='d29763;             
          'd3529 : value = 'h7454;    //value='d29780;             
          'd3530 : value = 'h7465;    //value='d29797;             
          'd3531 : value = 'h7476;    //value='d29814;             
          'd3532 : value = 'h7486;    //value='d29830;             
          'd3533 : value = 'h7497;    //value='d29847;             
          'd3534 : value = 'h74A8;    //value='d29864;             
          'd3535 : value = 'h74B9;    //value='d29881;             
          'd3536 : value = 'h74C9;    //value='d29897;             
          'd3537 : value = 'h74DA;    //value='d29914;             
          'd3538 : value = 'h74EB;    //value='d29931;             
          'd3539 : value = 'h74FC;    //value='d29948;             
          'd3540 : value = 'h750D;    //value='d29965;             
          'd3541 : value = 'h751E;    //value='d29982;             
          'd3542 : value = 'h752E;    //value='d29998;             
          'd3543 : value = 'h753F;    //value='d30015;             
          'd3544 : value = 'h7550;    //value='d30032;             
          'd3545 : value = 'h7561;    //value='d30049;             
          'd3546 : value = 'h7572;    //value='d30066;             
          'd3547 : value = 'h7583;    //value='d30083;             
          'd3548 : value = 'h7594;    //value='d30100;             
          'd3549 : value = 'h75A5;    //value='d30117;             
          'd3550 : value = 'h75B6;    //value='d30134;             
          'd3551 : value = 'h75C7;    //value='d30151;             
          'd3552 : value = 'h75D8;    //value='d30168;             
          'd3553 : value = 'h75E9;    //value='d30185;             
          'd3554 : value = 'h75FA;    //value='d30202;             
          'd3555 : value = 'h760A;    //value='d30218;             
          'd3556 : value = 'h761B;    //value='d30235;             
          'd3557 : value = 'h762C;    //value='d30252;             
          'd3558 : value = 'h763D;    //value='d30269;             
          'd3559 : value = 'h764F;    //value='d30287;             
          'd3560 : value = 'h7660;    //value='d30304;             
          'd3561 : value = 'h7671;    //value='d30321;             
          'd3562 : value = 'h7682;    //value='d30338;             
          'd3563 : value = 'h7693;    //value='d30355;             
          'd3564 : value = 'h76A4;    //value='d30372;             
          'd3565 : value = 'h76B5;    //value='d30389;             
          'd3566 : value = 'h76C6;    //value='d30406;             
          'd3567 : value = 'h76D7;    //value='d30423;             
          'd3568 : value = 'h76E8;    //value='d30440;             
          'd3569 : value = 'h76F9;    //value='d30457;             
          'd3570 : value = 'h770A;    //value='d30474;             
          'd3571 : value = 'h771C;    //value='d30492;             
          'd3572 : value = 'h772D;    //value='d30509;             
          'd3573 : value = 'h773E;    //value='d30526;             
          'd3574 : value = 'h774F;    //value='d30543;             
          'd3575 : value = 'h7760;    //value='d30560;             
          'd3576 : value = 'h7771;    //value='d30577;             
          'd3577 : value = 'h7783;    //value='d30595;             
          'd3578 : value = 'h7794;    //value='d30612;             
          'd3579 : value = 'h77A5;    //value='d30629;             
          'd3580 : value = 'h77B6;    //value='d30646;             
          'd3581 : value = 'h77C7;    //value='d30663;             
          'd3582 : value = 'h77D9;    //value='d30681;             
          'd3583 : value = 'h77EA;    //value='d30698;             
          'd3584 : value = 'h77FB;    //value='d30715;             
          'd3585 : value = 'h780C;    //value='d30732;             
          'd3586 : value = 'h781E;    //value='d30750;             
          'd3587 : value = 'h782F;    //value='d30767;             
          'd3588 : value = 'h7840;    //value='d30784;             
          'd3589 : value = 'h7852;    //value='d30802;             
          'd3590 : value = 'h7863;    //value='d30819;             
          'd3591 : value = 'h7874;    //value='d30836;             
          'd3592 : value = 'h7886;    //value='d30854;             
          'd3593 : value = 'h7897;    //value='d30871;             
          'd3594 : value = 'h78A8;    //value='d30888;             
          'd3595 : value = 'h78BA;    //value='d30906;             
          'd3596 : value = 'h78CB;    //value='d30923;             
          'd3597 : value = 'h78DC;    //value='d30940;             
          'd3598 : value = 'h78EE;    //value='d30958;             
          'd3599 : value = 'h78FF;    //value='d30975;             
          'd3600 : value = 'h7911;    //value='d30993;             
          'd3601 : value = 'h7922;    //value='d31010;             
          'd3602 : value = 'h7934;    //value='d31028;             
          'd3603 : value = 'h7945;    //value='d31045;             
          'd3604 : value = 'h7956;    //value='d31062;             
          'd3605 : value = 'h7968;    //value='d31080;             
          'd3606 : value = 'h7979;    //value='d31097;             
          'd3607 : value = 'h798B;    //value='d31115;             
          'd3608 : value = 'h799C;    //value='d31132;             
          'd3609 : value = 'h79AE;    //value='d31150;             
          'd3610 : value = 'h79BF;    //value='d31167;             
          'd3611 : value = 'h79D1;    //value='d31185;             
          'd3612 : value = 'h79E2;    //value='d31202;             
          'd3613 : value = 'h79F4;    //value='d31220;             
          'd3614 : value = 'h7A06;    //value='d31238;             
          'd3615 : value = 'h7A17;    //value='d31255;             
          'd3616 : value = 'h7A29;    //value='d31273;             
          'd3617 : value = 'h7A3A;    //value='d31290;             
          'd3618 : value = 'h7A4C;    //value='d31308;             
          'd3619 : value = 'h7A5D;    //value='d31325;             
          'd3620 : value = 'h7A6F;    //value='d31343;             
          'd3621 : value = 'h7A81;    //value='d31361;             
          'd3622 : value = 'h7A92;    //value='d31378;             
          'd3623 : value = 'h7AA4;    //value='d31396;             
          'd3624 : value = 'h7AB6;    //value='d31414;             
          'd3625 : value = 'h7AC7;    //value='d31431;             
          'd3626 : value = 'h7AD9;    //value='d31449;             
          'd3627 : value = 'h7AEB;    //value='d31467;             
          'd3628 : value = 'h7AFC;    //value='d31484;             
          'd3629 : value = 'h7B0E;    //value='d31502;             
          'd3630 : value = 'h7B20;    //value='d31520;             
          'd3631 : value = 'h7B32;    //value='d31538;             
          'd3632 : value = 'h7B43;    //value='d31555;             
          'd3633 : value = 'h7B55;    //value='d31573;             
          'd3634 : value = 'h7B67;    //value='d31591;             
          'd3635 : value = 'h7B79;    //value='d31609;             
          'd3636 : value = 'h7B8A;    //value='d31626;             
          'd3637 : value = 'h7B9C;    //value='d31644;             
          'd3638 : value = 'h7BAE;    //value='d31662;             
          'd3639 : value = 'h7BC0;    //value='d31680;             
          'd3640 : value = 'h7BD1;    //value='d31697;             
          'd3641 : value = 'h7BE3;    //value='d31715;             
          'd3642 : value = 'h7BF5;    //value='d31733;             
          'd3643 : value = 'h7C07;    //value='d31751;             
          'd3644 : value = 'h7C19;    //value='d31769;             
          'd3645 : value = 'h7C2B;    //value='d31787;             
          'd3646 : value = 'h7C3D;    //value='d31805;             
          'd3647 : value = 'h7C4E;    //value='d31822;             
          'd3648 : value = 'h7C60;    //value='d31840;             
          'd3649 : value = 'h7C72;    //value='d31858;             
          'd3650 : value = 'h7C84;    //value='d31876;             
          'd3651 : value = 'h7C96;    //value='d31894;             
          'd3652 : value = 'h7CA8;    //value='d31912;             
          'd3653 : value = 'h7CBA;    //value='d31930;             
          'd3654 : value = 'h7CCC;    //value='d31948;             
          'd3655 : value = 'h7CDE;    //value='d31966;             
          'd3656 : value = 'h7CF0;    //value='d31984;             
          'd3657 : value = 'h7D02;    //value='d32002;             
          'd3658 : value = 'h7D14;    //value='d32020;             
          'd3659 : value = 'h7D26;    //value='d32038;             
          'd3660 : value = 'h7D38;    //value='d32056;             
          'd3661 : value = 'h7D4A;    //value='d32074;             
          'd3662 : value = 'h7D5C;    //value='d32092;             
          'd3663 : value = 'h7D6E;    //value='d32110;             
          'd3664 : value = 'h7D80;    //value='d32128;             
          'd3665 : value = 'h7D92;    //value='d32146;             
          'd3666 : value = 'h7DA4;    //value='d32164;             
          'd3667 : value = 'h7DB6;    //value='d32182;             
          'd3668 : value = 'h7DC8;    //value='d32200;             
          'd3669 : value = 'h7DDA;    //value='d32218;             
          'd3670 : value = 'h7DED;    //value='d32237;             
          'd3671 : value = 'h7DFF;    //value='d32255;             
          'd3672 : value = 'h7E11;    //value='d32273;             
          'd3673 : value = 'h7E23;    //value='d32291;             
          'd3674 : value = 'h7E35;    //value='d32309;             
          'd3675 : value = 'h7E47;    //value='d32327;             
          'd3676 : value = 'h7E5A;    //value='d32346;             
          'd3677 : value = 'h7E6C;    //value='d32364;             
          'd3678 : value = 'h7E7E;    //value='d32382;             
          'd3679 : value = 'h7E90;    //value='d32400;             
          'd3680 : value = 'h7EA2;    //value='d32418;             
          'd3681 : value = 'h7EB5;    //value='d32437;             
          'd3682 : value = 'h7EC7;    //value='d32455;             
          'd3683 : value = 'h7ED9;    //value='d32473;             
          'd3684 : value = 'h7EEB;    //value='d32491;             
          'd3685 : value = 'h7EFE;    //value='d32510;             
          'd3686 : value = 'h7F10;    //value='d32528;             
          'd3687 : value = 'h7F22;    //value='d32546;             
          'd3688 : value = 'h7F34;    //value='d32564;             
          'd3689 : value = 'h7F47;    //value='d32583;             
          'd3690 : value = 'h7F59;    //value='d32601;             
          'd3691 : value = 'h7F6B;    //value='d32619;             
          'd3692 : value = 'h7F7E;    //value='d32638;             
          'd3693 : value = 'h7F90;    //value='d32656;             
          'd3694 : value = 'h7FA2;    //value='d32674;             
          'd3695 : value = 'h7FB5;    //value='d32693;             
          'd3696 : value = 'h7FC7;    //value='d32711;             
          'd3697 : value = 'h7FDA;    //value='d32730;             
          'd3698 : value = 'h7FEC;    //value='d32748;             
          'd3699 : value = 'h7FFE;    //value='d32766;             
          'd3700 : value = 'h8011;    //value='d32785;             
          'd3701 : value = 'h8023;    //value='d32803;             
          'd3702 : value = 'h8036;    //value='d32822;             
          'd3703 : value = 'h8048;    //value='d32840;             
          'd3704 : value = 'h805B;    //value='d32859;             
          'd3705 : value = 'h806D;    //value='d32877;             
          'd3706 : value = 'h8080;    //value='d32896;             
          'd3707 : value = 'h8092;    //value='d32914;             
          'd3708 : value = 'h80A5;    //value='d32933;             
          'd3709 : value = 'h80B7;    //value='d32951;             
          'd3710 : value = 'h80CA;    //value='d32970;             
          'd3711 : value = 'h80DC;    //value='d32988;             
          'd3712 : value = 'h80EF;    //value='d33007;             
          'd3713 : value = 'h8101;    //value='d33025;             
          'd3714 : value = 'h8114;    //value='d33044;             
          'd3715 : value = 'h8127;    //value='d33063;             
          'd3716 : value = 'h8139;    //value='d33081;             
          'd3717 : value = 'h814C;    //value='d33100;             
          'd3718 : value = 'h815E;    //value='d33118;             
          'd3719 : value = 'h8171;    //value='d33137;             
          'd3720 : value = 'h8184;    //value='d33156;             
          'd3721 : value = 'h8196;    //value='d33174;             
          'd3722 : value = 'h81A9;    //value='d33193;             
          'd3723 : value = 'h81BC;    //value='d33212;             
          'd3724 : value = 'h81CE;    //value='d33230;             
          'd3725 : value = 'h81E1;    //value='d33249;             
          'd3726 : value = 'h81F4;    //value='d33268;             
          'd3727 : value = 'h8206;    //value='d33286;             
          'd3728 : value = 'h8219;    //value='d33305;             
          'd3729 : value = 'h822C;    //value='d33324;             
          'd3730 : value = 'h823E;    //value='d33342;             
          'd3731 : value = 'h8251;    //value='d33361;             
          'd3732 : value = 'h8264;    //value='d33380;             
          'd3733 : value = 'h8277;    //value='d33399;             
          'd3734 : value = 'h828A;    //value='d33418;             
          'd3735 : value = 'h829C;    //value='d33436;             
          'd3736 : value = 'h82AF;    //value='d33455;             
          'd3737 : value = 'h82C2;    //value='d33474;             
          'd3738 : value = 'h82D5;    //value='d33493;             
          'd3739 : value = 'h82E8;    //value='d33512;             
          'd3740 : value = 'h82FA;    //value='d33530;             
          'd3741 : value = 'h830D;    //value='d33549;             
          'd3742 : value = 'h8320;    //value='d33568;             
          'd3743 : value = 'h8333;    //value='d33587;             
          'd3744 : value = 'h8346;    //value='d33606;             
          'd3745 : value = 'h8359;    //value='d33625;             
          'd3746 : value = 'h836C;    //value='d33644;             
          'd3747 : value = 'h837F;    //value='d33663;             
          'd3748 : value = 'h8392;    //value='d33682;             
          'd3749 : value = 'h83A5;    //value='d33701;             
          'd3750 : value = 'h83B7;    //value='d33719;             
          'd3751 : value = 'h83CA;    //value='d33738;             
          'd3752 : value = 'h83DD;    //value='d33757;             
          'd3753 : value = 'h83F0;    //value='d33776;             
          'd3754 : value = 'h8403;    //value='d33795;             
          'd3755 : value = 'h8416;    //value='d33814;             
          'd3756 : value = 'h8429;    //value='d33833;             
          'd3757 : value = 'h843C;    //value='d33852;             
          'd3758 : value = 'h844F;    //value='d33871;             
          'd3759 : value = 'h8463;    //value='d33891;             
          'd3760 : value = 'h8476;    //value='d33910;             
          'd3761 : value = 'h8489;    //value='d33929;             
          'd3762 : value = 'h849C;    //value='d33948;             
          'd3763 : value = 'h84AF;    //value='d33967;             
          'd3764 : value = 'h84C2;    //value='d33986;             
          'd3765 : value = 'h84D5;    //value='d34005;             
          'd3766 : value = 'h84E8;    //value='d34024;             
          'd3767 : value = 'h84FB;    //value='d34043;             
          'd3768 : value = 'h850E;    //value='d34062;             
          'd3769 : value = 'h8522;    //value='d34082;             
          'd3770 : value = 'h8535;    //value='d34101;             
          'd3771 : value = 'h8548;    //value='d34120;             
          'd3772 : value = 'h855B;    //value='d34139;             
          'd3773 : value = 'h856E;    //value='d34158;             
          'd3774 : value = 'h8582;    //value='d34178;             
          'd3775 : value = 'h8595;    //value='d34197;             
          'd3776 : value = 'h85A8;    //value='d34216;             
          'd3777 : value = 'h85BB;    //value='d34235;             
          'd3778 : value = 'h85CE;    //value='d34254;             
          'd3779 : value = 'h85E2;    //value='d34274;             
          'd3780 : value = 'h85F5;    //value='d34293;             
          'd3781 : value = 'h8608;    //value='d34312;             
          'd3782 : value = 'h861C;    //value='d34332;             
          'd3783 : value = 'h862F;    //value='d34351;             
          'd3784 : value = 'h8642;    //value='d34370;             
          'd3785 : value = 'h8656;    //value='d34390;             
          'd3786 : value = 'h8669;    //value='d34409;             
          'd3787 : value = 'h867C;    //value='d34428;             
          'd3788 : value = 'h8690;    //value='d34448;             
          'd3789 : value = 'h86A3;    //value='d34467;             
          'd3790 : value = 'h86B6;    //value='d34486;             
          'd3791 : value = 'h86CA;    //value='d34506;             
          'd3792 : value = 'h86DD;    //value='d34525;             
          'd3793 : value = 'h86F1;    //value='d34545;             
          'd3794 : value = 'h8704;    //value='d34564;             
          'd3795 : value = 'h8717;    //value='d34583;             
          'd3796 : value = 'h872B;    //value='d34603;             
          'd3797 : value = 'h873E;    //value='d34622;             
          'd3798 : value = 'h8752;    //value='d34642;             
          'd3799 : value = 'h8765;    //value='d34661;             
          'd3800 : value = 'h8779;    //value='d34681;             
          'd3801 : value = 'h878C;    //value='d34700;             
          'd3802 : value = 'h87A0;    //value='d34720;             
          'd3803 : value = 'h87B3;    //value='d34739;             
          'd3804 : value = 'h87C7;    //value='d34759;             
          'd3805 : value = 'h87DA;    //value='d34778;             
          'd3806 : value = 'h87EE;    //value='d34798;             
          'd3807 : value = 'h8801;    //value='d34817;             
          'd3808 : value = 'h8815;    //value='d34837;             
          'd3809 : value = 'h8829;    //value='d34857;             
          'd3810 : value = 'h883C;    //value='d34876;             
          'd3811 : value = 'h8850;    //value='d34896;             
          'd3812 : value = 'h8863;    //value='d34915;             
          'd3813 : value = 'h8877;    //value='d34935;             
          'd3814 : value = 'h888B;    //value='d34955;             
          'd3815 : value = 'h889E;    //value='d34974;             
          'd3816 : value = 'h88B2;    //value='d34994;             
          'd3817 : value = 'h88C6;    //value='d35014;             
          'd3818 : value = 'h88D9;    //value='d35033;             
          'd3819 : value = 'h88ED;    //value='d35053;             
          'd3820 : value = 'h8901;    //value='d35073;             
          'd3821 : value = 'h8915;    //value='d35093;             
          'd3822 : value = 'h8928;    //value='d35112;             
          'd3823 : value = 'h893C;    //value='d35132;             
          'd3824 : value = 'h8950;    //value='d35152;             
          'd3825 : value = 'h8964;    //value='d35172;             
          'd3826 : value = 'h8977;    //value='d35191;             
          'd3827 : value = 'h898B;    //value='d35211;             
          'd3828 : value = 'h899F;    //value='d35231;             
          'd3829 : value = 'h89B3;    //value='d35251;             
          'd3830 : value = 'h89C7;    //value='d35271;             
          'd3831 : value = 'h89DA;    //value='d35290;             
          'd3832 : value = 'h89EE;    //value='d35310;             
          'd3833 : value = 'h8A02;    //value='d35330;             
          'd3834 : value = 'h8A16;    //value='d35350;             
          'd3835 : value = 'h8A2A;    //value='d35370;             
          'd3836 : value = 'h8A3E;    //value='d35390;             
          'd3837 : value = 'h8A52;    //value='d35410;             
          'd3838 : value = 'h8A66;    //value='d35430;             
          'd3839 : value = 'h8A79;    //value='d35449;             
          'd3840 : value = 'h8A8D;    //value='d35469;             
          'd3841 : value = 'h8AA1;    //value='d35489;             
          'd3842 : value = 'h8AB5;    //value='d35509;             
          'd3843 : value = 'h8AC9;    //value='d35529;             
          'd3844 : value = 'h8ADD;    //value='d35549;             
          'd3845 : value = 'h8AF1;    //value='d35569;             
          'd3846 : value = 'h8B05;    //value='d35589;             
          'd3847 : value = 'h8B19;    //value='d35609;             
          'd3848 : value = 'h8B2D;    //value='d35629;             
          'd3849 : value = 'h8B41;    //value='d35649;             
          'd3850 : value = 'h8B55;    //value='d35669;             
          'd3851 : value = 'h8B69;    //value='d35689;             
          'd3852 : value = 'h8B7D;    //value='d35709;             
          'd3853 : value = 'h8B92;    //value='d35730;             
          'd3854 : value = 'h8BA6;    //value='d35750;             
          'd3855 : value = 'h8BBA;    //value='d35770;             
          'd3856 : value = 'h8BCE;    //value='d35790;             
          'd3857 : value = 'h8BE2;    //value='d35810;             
          'd3858 : value = 'h8BF6;    //value='d35830;             
          'd3859 : value = 'h8C0A;    //value='d35850;             
          'd3860 : value = 'h8C1E;    //value='d35870;             
          'd3861 : value = 'h8C33;    //value='d35891;             
          'd3862 : value = 'h8C47;    //value='d35911;             
          'd3863 : value = 'h8C5B;    //value='d35931;             
          'd3864 : value = 'h8C6F;    //value='d35951;             
          'd3865 : value = 'h8C83;    //value='d35971;             
          'd3866 : value = 'h8C98;    //value='d35992;             
          'd3867 : value = 'h8CAC;    //value='d36012;             
          'd3868 : value = 'h8CC0;    //value='d36032;             
          'd3869 : value = 'h8CD4;    //value='d36052;             
          'd3870 : value = 'h8CE9;    //value='d36073;             
          'd3871 : value = 'h8CFD;    //value='d36093;             
          'd3872 : value = 'h8D11;    //value='d36113;             
          'd3873 : value = 'h8D26;    //value='d36134;             
          'd3874 : value = 'h8D3A;    //value='d36154;             
          'd3875 : value = 'h8D4E;    //value='d36174;             
          'd3876 : value = 'h8D63;    //value='d36195;             
          'd3877 : value = 'h8D77;    //value='d36215;             
          'd3878 : value = 'h8D8B;    //value='d36235;             
          'd3879 : value = 'h8DA0;    //value='d36256;             
          'd3880 : value = 'h8DB4;    //value='d36276;             
          'd3881 : value = 'h8DC8;    //value='d36296;             
          'd3882 : value = 'h8DDD;    //value='d36317;             
          'd3883 : value = 'h8DF1;    //value='d36337;             
          'd3884 : value = 'h8E06;    //value='d36358;             
          'd3885 : value = 'h8E1A;    //value='d36378;             
          'd3886 : value = 'h8E2F;    //value='d36399;             
          'd3887 : value = 'h8E43;    //value='d36419;             
          'd3888 : value = 'h8E58;    //value='d36440;             
          'd3889 : value = 'h8E6C;    //value='d36460;             
          'd3890 : value = 'h8E81;    //value='d36481;             
          'd3891 : value = 'h8E95;    //value='d36501;             
          'd3892 : value = 'h8EAA;    //value='d36522;             
          'd3893 : value = 'h8EBE;    //value='d36542;             
          'd3894 : value = 'h8ED3;    //value='d36563;             
          'd3895 : value = 'h8EE7;    //value='d36583;             
          'd3896 : value = 'h8EFC;    //value='d36604;             
          'd3897 : value = 'h8F10;    //value='d36624;             
          'd3898 : value = 'h8F25;    //value='d36645;             
          'd3899 : value = 'h8F3A;    //value='d36666;             
          'd3900 : value = 'h8F4E;    //value='d36686;             
          'd3901 : value = 'h8F63;    //value='d36707;             
          'd3902 : value = 'h8F77;    //value='d36727;             
          'd3903 : value = 'h8F8C;    //value='d36748;             
          'd3904 : value = 'h8FA1;    //value='d36769;             
          'd3905 : value = 'h8FB5;    //value='d36789;             
          'd3906 : value = 'h8FCA;    //value='d36810;             
          'd3907 : value = 'h8FDF;    //value='d36831;             
          'd3908 : value = 'h8FF4;    //value='d36852;             
          'd3909 : value = 'h9008;    //value='d36872;             
          'd3910 : value = 'h901D;    //value='d36893;             
          'd3911 : value = 'h9032;    //value='d36914;             
          'd3912 : value = 'h9046;    //value='d36934;             
          'd3913 : value = 'h905B;    //value='d36955;             
          'd3914 : value = 'h9070;    //value='d36976;             
          'd3915 : value = 'h9085;    //value='d36997;             
          'd3916 : value = 'h909A;    //value='d37018;             
          'd3917 : value = 'h90AE;    //value='d37038;             
          'd3918 : value = 'h90C3;    //value='d37059;             
          'd3919 : value = 'h90D8;    //value='d37080;             
          'd3920 : value = 'h90ED;    //value='d37101;             
          'd3921 : value = 'h9102;    //value='d37122;             
          'd3922 : value = 'h9117;    //value='d37143;             
          'd3923 : value = 'h912C;    //value='d37164;             
          'd3924 : value = 'h9140;    //value='d37184;             
          'd3925 : value = 'h9155;    //value='d37205;             
          'd3926 : value = 'h916A;    //value='d37226;             
          'd3927 : value = 'h917F;    //value='d37247;             
          'd3928 : value = 'h9194;    //value='d37268;             
          'd3929 : value = 'h91A9;    //value='d37289;             
          'd3930 : value = 'h91BE;    //value='d37310;             
          'd3931 : value = 'h91D3;    //value='d37331;             
          'd3932 : value = 'h91E8;    //value='d37352;             
          'd3933 : value = 'h91FD;    //value='d37373;             
          'd3934 : value = 'h9212;    //value='d37394;             
          'd3935 : value = 'h9227;    //value='d37415;             
          'd3936 : value = 'h923C;    //value='d37436;             
          'd3937 : value = 'h9251;    //value='d37457;             
          'd3938 : value = 'h9266;    //value='d37478;             
          'd3939 : value = 'h927B;    //value='d37499;             
          'd3940 : value = 'h9290;    //value='d37520;             
          'd3941 : value = 'h92A6;    //value='d37542;             
          'd3942 : value = 'h92BB;    //value='d37563;             
          'd3943 : value = 'h92D0;    //value='d37584;             
          'd3944 : value = 'h92E5;    //value='d37605;             
          'd3945 : value = 'h92FA;    //value='d37626;             
          'd3946 : value = 'h930F;    //value='d37647;             
          'd3947 : value = 'h9324;    //value='d37668;             
          'd3948 : value = 'h933A;    //value='d37690;             
          'd3949 : value = 'h934F;    //value='d37711;             
          'd3950 : value = 'h9364;    //value='d37732;             
          'd3951 : value = 'h9379;    //value='d37753;             
          'd3952 : value = 'h938E;    //value='d37774;             
          'd3953 : value = 'h93A4;    //value='d37796;             
          'd3954 : value = 'h93B9;    //value='d37817;             
          'd3955 : value = 'h93CE;    //value='d37838;             
          'd3956 : value = 'h93E3;    //value='d37859;             
          'd3957 : value = 'h93F9;    //value='d37881;             
          'd3958 : value = 'h940E;    //value='d37902;             
          'd3959 : value = 'h9423;    //value='d37923;             
          'd3960 : value = 'h9439;    //value='d37945;             
          'd3961 : value = 'h944E;    //value='d37966;             
          'd3962 : value = 'h9463;    //value='d37987;             
          'd3963 : value = 'h9479;    //value='d38009;             
          'd3964 : value = 'h948E;    //value='d38030;             
          'd3965 : value = 'h94A4;    //value='d38052;             
          'd3966 : value = 'h94B9;    //value='d38073;             
          'd3967 : value = 'h94CE;    //value='d38094;             
          'd3968 : value = 'h94E4;    //value='d38116;             
          'd3969 : value = 'h94F9;    //value='d38137;             
          'd3970 : value = 'h950F;    //value='d38159;             
          'd3971 : value = 'h9524;    //value='d38180;             
          'd3972 : value = 'h953A;    //value='d38202;             
          'd3973 : value = 'h954F;    //value='d38223;             
          'd3974 : value = 'h9565;    //value='d38245;             
          'd3975 : value = 'h957A;    //value='d38266;             
          'd3976 : value = 'h9590;    //value='d38288;             
          'd3977 : value = 'h95A5;    //value='d38309;             
          'd3978 : value = 'h95BB;    //value='d38331;             
          'd3979 : value = 'h95D0;    //value='d38352;             
          'd3980 : value = 'h95E6;    //value='d38374;             
          'd3981 : value = 'h95FB;    //value='d38395;             
          'd3982 : value = 'h9611;    //value='d38417;             
          'd3983 : value = 'h9626;    //value='d38438;             
          'd3984 : value = 'h963C;    //value='d38460;             
          'd3985 : value = 'h9652;    //value='d38482;             
          'd3986 : value = 'h9667;    //value='d38503;             
          'd3987 : value = 'h967D;    //value='d38525;             
          'd3988 : value = 'h9693;    //value='d38547;             
          'd3989 : value = 'h96A8;    //value='d38568;             
          'd3990 : value = 'h96BE;    //value='d38590;             
          'd3991 : value = 'h96D4;    //value='d38612;             
          'd3992 : value = 'h96E9;    //value='d38633;             
          'd3993 : value = 'h96FF;    //value='d38655;             
          'd3994 : value = 'h9715;    //value='d38677;             
          'd3995 : value = 'h972B;    //value='d38699;             
          'd3996 : value = 'h9740;    //value='d38720;             
          'd3997 : value = 'h9756;    //value='d38742;             
          'd3998 : value = 'h976C;    //value='d38764;             
          'd3999 : value = 'h9782;    //value='d38786;             
          'd4000 : value = 'h9798;    //value='d38808;             
          'd4001 : value = 'h97AD;    //value='d38829;             
          'd4002 : value = 'h97C3;    //value='d38851;             
          'd4003 : value = 'h97D9;    //value='d38873;             
          'd4004 : value = 'h97EF;    //value='d38895;             
          'd4005 : value = 'h9805;    //value='d38917;             
          'd4006 : value = 'h981B;    //value='d38939;             
          'd4007 : value = 'h9831;    //value='d38961;             
          'd4008 : value = 'h9847;    //value='d38983;             
          'd4009 : value = 'h985C;    //value='d39004;             
          'd4010 : value = 'h9872;    //value='d39026;             
          'd4011 : value = 'h9888;    //value='d39048;             
          'd4012 : value = 'h989E;    //value='d39070;             
          'd4013 : value = 'h98B4;    //value='d39092;             
          'd4014 : value = 'h98CA;    //value='d39114;             
          'd4015 : value = 'h98E0;    //value='d39136;             
          'd4016 : value = 'h98F6;    //value='d39158;             
          'd4017 : value = 'h990C;    //value='d39180;             
          'd4018 : value = 'h9922;    //value='d39202;             
          'd4019 : value = 'h9938;    //value='d39224;             
          'd4020 : value = 'h994E;    //value='d39246;             
          'd4021 : value = 'h9964;    //value='d39268;             
          'd4022 : value = 'h997B;    //value='d39291;             
          'd4023 : value = 'h9991;    //value='d39313;             
          'd4024 : value = 'h99A7;    //value='d39335;             
          'd4025 : value = 'h99BD;    //value='d39357;             
          'd4026 : value = 'h99D3;    //value='d39379;             
          'd4027 : value = 'h99E9;    //value='d39401;             
          'd4028 : value = 'h99FF;    //value='d39423;             
          'd4029 : value = 'h9A15;    //value='d39445;             
          'd4030 : value = 'h9A2C;    //value='d39468;             
          'd4031 : value = 'h9A42;    //value='d39490;             
          'd4032 : value = 'h9A58;    //value='d39512;             
          'd4033 : value = 'h9A6E;    //value='d39534;             
          'd4034 : value = 'h9A84;    //value='d39556;             
          'd4035 : value = 'h9A9B;    //value='d39579;             
          'd4036 : value = 'h9AB1;    //value='d39601;             
          'd4037 : value = 'h9AC7;    //value='d39623;             
          'd4038 : value = 'h9ADE;    //value='d39646;             
          'd4039 : value = 'h9AF4;    //value='d39668;             
          'd4040 : value = 'h9B0A;    //value='d39690;             
          'd4041 : value = 'h9B20;    //value='d39712;             
          'd4042 : value = 'h9B37;    //value='d39735;             
          'd4043 : value = 'h9B4D;    //value='d39757;             
          'd4044 : value = 'h9B63;    //value='d39779;             
          'd4045 : value = 'h9B7A;    //value='d39802;             
          'd4046 : value = 'h9B90;    //value='d39824;             
          'd4047 : value = 'h9BA7;    //value='d39847;             
          'd4048 : value = 'h9BBD;    //value='d39869;             
          'd4049 : value = 'h9BD3;    //value='d39891;             
          'd4050 : value = 'h9BEA;    //value='d39914;             
          'd4051 : value = 'h9C00;    //value='d39936;             
          'd4052 : value = 'h9C17;    //value='d39959;             
          'd4053 : value = 'h9C2D;    //value='d39981;             
          'd4054 : value = 'h9C44;    //value='d40004;             
          'd4055 : value = 'h9C5A;    //value='d40026;             
          'd4056 : value = 'h9C71;    //value='d40049;             
          'd4057 : value = 'h9C87;    //value='d40071;             
          'd4058 : value = 'h9C9E;    //value='d40094;             
          'd4059 : value = 'h9CB4;    //value='d40116;             
          'd4060 : value = 'h9CCB;    //value='d40139;             
          'd4061 : value = 'h9CE1;    //value='d40161;             
          'd4062 : value = 'h9CF8;    //value='d40184;             
          'd4063 : value = 'h9D0F;    //value='d40207;             
          'd4064 : value = 'h9D25;    //value='d40229;             
          'd4065 : value = 'h9D3C;    //value='d40252;             
          'd4066 : value = 'h9D53;    //value='d40275;             
          'd4067 : value = 'h9D69;    //value='d40297;             
          'd4068 : value = 'h9D80;    //value='d40320;             
          'd4069 : value = 'h9D96;    //value='d40342;             
          'd4070 : value = 'h9DAD;    //value='d40365;             
          'd4071 : value = 'h9DC4;    //value='d40388;             
          'd4072 : value = 'h9DDB;    //value='d40411;             
          'd4073 : value = 'h9DF1;    //value='d40433;             
          'd4074 : value = 'h9E08;    //value='d40456;             
          'd4075 : value = 'h9E1F;    //value='d40479;             
          'd4076 : value = 'h9E36;    //value='d40502;             
          'd4077 : value = 'h9E4C;    //value='d40524;             
          'd4078 : value = 'h9E63;    //value='d40547;             
          'd4079 : value = 'h9E7A;    //value='d40570;             
          'd4080 : value = 'h9E91;    //value='d40593;             
          'd4081 : value = 'h9EA8;    //value='d40616;             
          'd4082 : value = 'h9EBE;    //value='d40638;             
          'd4083 : value = 'h9ED5;    //value='d40661;             
          'd4084 : value = 'h9EEC;    //value='d40684;             
          'd4085 : value = 'h9F03;    //value='d40707;             
          'd4086 : value = 'h9F1A;    //value='d40730;             
          'd4087 : value = 'h9F31;    //value='d40753;             
          'd4088 : value = 'h9F48;    //value='d40776;             
          'd4089 : value = 'h9F5F;    //value='d40799;             
          'd4090 : value = 'h9F76;    //value='d40822;             
          'd4091 : value = 'h9F8D;    //value='d40845;             
          'd4092 : value = 'h9FA4;    //value='d40868;             
          'd4093 : value = 'h9FBA;    //value='d40890;             
          'd4094 : value = 'h9FD1;    //value='d40913;             
          'd4095 : value = 'h9FE8;    //value='d40936;             
endcase   
end   


endmodule   
