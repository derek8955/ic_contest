

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO IOTDF 
  PIN iot_in[7] 
    ANTENNAPARTIALMETALAREA 8.044 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.154 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 13.112 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.032 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 31.651 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 111.059 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2756 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 254.016 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 895.189 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.78645 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 9.224 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 32.564 LAYER METAL5 ;
    ANTENNAGATEAREA 0.8411 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 264.983 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 933.905 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.36597 LAYER VIA56 ;
  END iot_in[7]
  PIN iot_in[6] 
    ANTENNAPARTIALMETALAREA 21.328 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 74.648 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 15.658 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.943 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 376.235 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 1321.94 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.52448 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 21.043 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 73.9305 LAYER METAL4 ;
    ANTENNAGATEAREA 0.4043 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 428.283 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1504.8 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.61377 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 17.262 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 60.557 LAYER METAL5 ;
    ANTENNAGATEAREA 0.8502 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 448.587 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1576.03 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.45761 LAYER VIA56 ;
  END iot_in[6]
  PIN iot_in[5] 
    ANTENNAPARTIALMETALAREA 18.13 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 63.455 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 17.328 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.068 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1287 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 211.783 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 746.357 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 3.92696 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 22.016 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 77.476 LAYER METAL4 ;
    ANTENNAGATEAREA 0.3614 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 272.702 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 960.734 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 4.02685 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 12.734 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 44.709 LAYER METAL5 ;
    ANTENNAGATEAREA 0.8502 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 287.68 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1013.32 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 4.02685 LAYER VIA56 ;
  END iot_in[5]
  PIN iot_in[4] 
    ANTENNAPARTIALMETALAREA 12.39 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 43.365 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 6.12 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.56 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 19.894 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 70.189 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2665 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 231.405 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 817.135 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 3.63689 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 34.306 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 120.491 LAYER METAL5 ;
    ANTENNAGATEAREA 0.8502 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 271.756 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 958.856 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.63689 LAYER VIA56 ;
  END iot_in[4]
  PIN iot_in[3] 
    ANTENNAPARTIALMETALAREA 10.012 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.042 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 6.12 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.56 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 19.553 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 68.8555 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5746 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 173.738 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 612.296 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.5873 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 6.57 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.135 LAYER METAL5 ;
    ANTENNAGATEAREA 0.8502 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 189.941 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 669.3 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.65546 LAYER VIA56 ;
  END iot_in[3]
  PIN iot_in[2] 
    ANTENNAPARTIALMETALAREA 3.944 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.804 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.278 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.613 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 41.954 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 147.539 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8502 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 192.097 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 676.538 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.91744 LAYER VIA45 ;
  END iot_in[2]
  PIN iot_in[1] 
    ANTENNAPARTIALMETALAREA 9.684 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.894 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.798 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.933 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 30.3 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 106.89 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7462 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 185.699 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 656.188 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 3.41435 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 9.718 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 34.153 LAYER METAL5 ;
    ANTENNAGATEAREA 0.8749 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 199.557 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 706.99 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.41435 LAYER VIA56 ;
  END iot_in[1]
  PIN iot_in[0] 
    ANTENNAPARTIALMETALAREA 4.19 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.665 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.702 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.597 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 35.596 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 125.006 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4563 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 260.085 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 914.086 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.92649 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 13.858 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 48.643 LAYER METAL5 ;
    ANTENNAGATEAREA 0.8502 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 276.385 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 971.3 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.08547 LAYER VIA56 ;
  END iot_in[0]
  PIN fn_sel[2] 
    ANTENNAPARTIALMETALAREA 9.284 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.494 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 10.362 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.407 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 24.82 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 87.01 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6292 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 54.3104 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 190.399 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.751605 LAYER VIA45 ;
  END fn_sel[2]
  PIN fn_sel[1] 
    ANTENNAPARTIALMETALAREA 10.094 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.329 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 13.459 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.2465 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 23.14 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 81.13 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5954 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 47.7279 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 168.66 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.52217 LAYER VIA45 ;
  END fn_sel[1]
  PIN fn_sel[0] 
    ANTENNAPARTIALMETALAREA 8.044 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.154 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 12.1 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.49 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 25.57 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 89.635 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8411 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 40.9234 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 144.245 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.660014 LAYER VIA45 ;
  END fn_sel[0]
  PIN iot_out[127] 
    ANTENNAPARTIALMETALAREA 9.356 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.746 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 9.35 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.865 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 21.06 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 73.85 LAYER METAL4 ;
  END iot_out[127]
  PIN iot_out[126] 
    ANTENNAPARTIALMETALAREA 9.858 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.503 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.382 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.477 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 17.624 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 61.824 LAYER METAL4 ;
  END iot_out[126]
  PIN iot_out[125] 
    ANTENNAPARTIALMETALAREA 9.93 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.755 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 7.326 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.781 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 20.946 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 73.451 LAYER METAL4 ;
  END iot_out[125]
  PIN iot_out[124] 
    ANTENNAPARTIALMETALAREA 3.534 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.369 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 7.878 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.713 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 27.138 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 95.123 LAYER METAL4 ;
  END iot_out[124]
  PIN iot_out[123] 
    ANTENNAPARTIALMETALAREA 9.284 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.494 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 7.142 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.137 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 21.316 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 74.746 LAYER METAL4 ;
  END iot_out[123]
  PIN iot_out[122] 
    ANTENNAPARTIALMETALAREA 9.438 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.033 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 6.478 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.813 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 21.622 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 75.817 LAYER METAL4 ;
  END iot_out[122]
  PIN iot_out[121] 
    ANTENNAPARTIALMETALAREA 8.044 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.154 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 5.384 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.984 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 22.442 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 78.687 LAYER METAL4 ;
  END iot_out[121]
  PIN iot_out[120] 
    ANTENNAPARTIALMETALAREA 10.278 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.973 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 8.226 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.931 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 19.994 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 70.119 LAYER METAL4 ;
  END iot_out[120]
  PIN iot_out[119] 
    ANTENNAPARTIALMETALAREA 8.618 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.163 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 7.694 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.069 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 22.648 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 79.408 LAYER METAL4 ;
  END iot_out[119]
  PIN iot_out[118] 
    ANTENNAPARTIALMETALAREA 8.382 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.337 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 6.957 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.4895 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 22.874 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 80.199 LAYER METAL4 ;
  END iot_out[118]
  PIN iot_out[117] 
    ANTENNAPARTIALMETALAREA 9.274 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.459 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 5.936 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.916 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 23.13 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 81.095 LAYER METAL4 ;
  END iot_out[117]
  PIN iot_out[116] 
    ANTENNAPARTIALMETALAREA 9.848 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.468 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.708 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.118 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 24.636 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 86.366 LAYER METAL4 ;
  END iot_out[116]
  PIN iot_out[115] 
    ANTENNAPARTIALMETALAREA 3.78 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.23 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.886 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.241 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 31.176 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 109.256 LAYER METAL4 ;
  END iot_out[115]
  PIN iot_out[114] 
    ANTENNAPARTIALMETALAREA 10.996 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.486 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.254 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.529 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 24.042 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 84.287 LAYER METAL4 ;
  END iot_out[114]
  PIN iot_out[113] 
    ANTENNAPARTIALMETALAREA 14.132 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.462 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.518 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.953 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 24.482 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 85.827 LAYER METAL4 ;
  END iot_out[113]
  PIN iot_out[112] 
    ANTENNAPARTIALMETALAREA 17.494 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.229 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.987 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 20.24 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 70.98 LAYER METAL4 ;
  END iot_out[112]
  PIN iot_out[111] 
    ANTENNAPARTIALMETALAREA 33.71 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 117.985 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.648 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.408 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 6.29 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.155 LAYER METAL4 ;
  END iot_out[111]
  PIN iot_out[110] 
    ANTENNAPARTIALMETALAREA 41.09 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 143.815 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 7.02 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.71 LAYER METAL3 ;
  END iot_out[110]
  PIN iot_out[109] 
    ANTENNAPARTIALMETALAREA 43.3 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 151.69 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 6.018 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.203 LAYER METAL3 ;
  END iot_out[109]
  PIN iot_out[108] 
    ANTENNAPARTIALMETALAREA 43.826 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.99 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.605 LAYER METAL3 ;
  END iot_out[108]
  PIN iot_out[107] 
    ANTENNAPARTIALMETALAREA 39.807 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 139.325 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 12.686 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 44.541 LAYER METAL4 ;
  END iot_out[107]
  PIN iot_out[106] 
    ANTENNAPARTIALMETALAREA 35.76 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 125.16 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 11.896 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.776 LAYER METAL4 ;
  END iot_out[106]
  PIN iot_out[105] 
    ANTENNAPARTIALMETALAREA 36.22 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 126.77 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 9.99 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 35.105 LAYER METAL4 ;
  END iot_out[105]
  PIN iot_out[104] 
    ANTENNAPARTIALMETALAREA 37.576 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 131.516 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 7.94 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.93 LAYER METAL4 ;
  END iot_out[104]
  PIN iot_out[103] 
    ANTENNAPARTIALMETALAREA 36.68 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 128.38 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 6.576 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 23.156 LAYER METAL4 ;
  END iot_out[103]
  PIN iot_out[102] 
    ANTENNAPARTIALMETALAREA 34.84 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 121.94 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 4.568 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.128 LAYER METAL4 ;
  END iot_out[102]
  PIN iot_out[101] 
    ANTENNAPARTIALMETALAREA 34.544 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 120.904 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.436 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.666 LAYER METAL4 ;
  END iot_out[101]
  PIN iot_out[100] 
    ANTENNAPARTIALMETALAREA 32.674 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 114.359 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.42 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.11 LAYER METAL4 ;
  END iot_out[100]
  PIN iot_out[99] 
    ANTENNAPARTIALMETALAREA 32.808 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 114.828 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 1.616 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.796 LAYER METAL4 ;
  END iot_out[99]
  PIN iot_out[98] 
    ANTENNAPARTIALMETALAREA 7.792 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.272 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.714 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.639 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 21.77 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 76.335 LAYER METAL5 ;
  END iot_out[98]
  PIN iot_out[97] 
    ANTENNAPARTIALMETALAREA 7.516 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.306 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.491 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 17.722 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 62.167 LAYER METAL5 ;
  END iot_out[97]
  PIN iot_out[96] 
    ANTENNAPARTIALMETALAREA 7.332 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.662 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.122 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.067 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 14.41 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 50.575 LAYER METAL5 ;
  END iot_out[96]
  PIN iot_out[95] 
    ANTENNAPARTIALMETALAREA 10.022 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.077 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 17.538 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 61.523 LAYER METAL5 ;
  END iot_out[95]
  PIN iot_out[94] 
    ANTENNAPARTIALMETALAREA 0.198 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.693 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.304 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 27.75 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 97.265 LAYER METAL5 ;
  END iot_out[94]
  PIN iot_out[93] 
    ANTENNAPARTIALMETALAREA 7.332 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.662 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.796 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.926 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 15.422 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 54.117 LAYER METAL5 ;
  END iot_out[93]
  PIN iot_out[92] 
    ANTENNAPARTIALMETALAREA 9.336 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.676 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 15.054 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 52.829 LAYER METAL5 ;
  END iot_out[92]
  PIN iot_out[91] 
    ANTENNAPARTIALMETALAREA 8.518 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.813 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.206 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.361 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 15.514 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 54.439 LAYER METAL5 ;
  END iot_out[91]
  PIN iot_out[90] 
    ANTENNAPARTIALMETALAREA 9.52 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.32 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 5.172 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.242 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 13.398 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 47.033 LAYER METAL5 ;
  END iot_out[90]
  PIN iot_out[89] 
    ANTENNAPARTIALMETALAREA 8.988 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.458 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 10.882 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.227 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 11.834 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 41.559 LAYER METAL5 ;
  END iot_out[89]
  PIN iot_out[88] 
    ANTENNAPARTIALMETALAREA 8.702 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.457 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 16.324 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 57.274 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 10.638 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 37.373 LAYER METAL5 ;
  END iot_out[88]
  PIN iot_out[87] 
    ANTENNAPARTIALMETALAREA 9.172 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.102 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 10.178 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 35.763 LAYER METAL5 ;
  END iot_out[87]
  PIN iot_out[86] 
    ANTENNAPARTIALMETALAREA 7.65 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.775 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.714 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.639 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.5916 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 9.626 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 33.831 LAYER METAL5 ;
  END iot_out[86]
  PIN iot_out[85] 
    ANTENNAPARTIALMETALAREA 9.264 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 5.946 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.951 LAYER METAL5 ;
  END iot_out[85]
  PIN iot_out[84] 
    ANTENNADIFFAREA 0.233 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.922 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.867 LAYER METAL3 ;
  END iot_out[84]
  PIN iot_out[83] 
    ANTENNAPARTIALMETALAREA 14.682 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.387 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 21.542 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 75.537 LAYER METAL4 ;
  END iot_out[83]
  PIN iot_out[82] 
    ANTENNAPARTIALMETALAREA 12.474 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.659 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 23.108 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 81.018 LAYER METAL4 ;
  END iot_out[82]
  PIN iot_out[81] 
    ANTENNADIFFAREA 0.233 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.34 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.83 LAYER METAL3 ;
  END iot_out[81]
  PIN iot_out[80] 
    ANTENNADIFFAREA 0.233 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.41 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.575 LAYER METAL3 ;
  END iot_out[80]
  PIN iot_out[79] 
    ANTENNAPARTIALMETALAREA 11.472 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.152 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 23.858 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 83.643 LAYER METAL4 ;
  END iot_out[79]
  PIN iot_out[78] 
    ANTENNAPARTIALMETALAREA 11.84 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.44 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 24.462 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 85.757 LAYER METAL4 ;
  END iot_out[78]
  PIN iot_out[77] 
    ANTENNAPARTIALMETALAREA 12.944 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.304 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 25.59 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 89.705 LAYER METAL4 ;
  END iot_out[77]
  PIN iot_out[76] 
    ANTENNAPARTIALMETALAREA 12.208 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.728 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 26.388 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 92.498 LAYER METAL4 ;
  END iot_out[76]
  PIN iot_out[75] 
    ANTENNADIFFAREA 0.233 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.57 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.135 LAYER METAL3 ;
  END iot_out[75]
  PIN iot_out[74] 
    ANTENNAPARTIALMETALAREA 13.864 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.524 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 26.882 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 94.227 LAYER METAL4 ;
  END iot_out[74]
  PIN iot_out[73] 
    ANTENNADIFFAREA 0.233 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.89 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.255 LAYER METAL3 ;
  END iot_out[73]
  PIN iot_out[72] 
    ANTENNAPARTIALMETALAREA 11.775 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.2125 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 28.758 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 100.793 LAYER METAL4 ;
  END iot_out[72]
  PIN iot_out[71] 
    ANTENNAPARTIALMETALAREA 23.818 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 83.363 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 16.496 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.876 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 4.814 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.989 LAYER METAL4 ;
  END iot_out[71]
  PIN iot_out[70] 
    ANTENNAPARTIALMETALAREA 9.776 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.216 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 15.79 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.405 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 17.974 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 63.049 LAYER METAL4 ;
  END iot_out[70]
  PIN iot_out[69] 
    ANTENNAPARTIALMETALAREA 7.224 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.284 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 12.928 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.388 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 18.732 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 65.702 LAYER METAL4 ;
  END iot_out[69]
  PIN iot_out[68] 
    ANTENNAPARTIALMETALAREA 8.044 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.154 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 8.236 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.966 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 16.324 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 57.274 LAYER METAL4 ;
  END iot_out[68]
  PIN iot_out[67] 
    ANTENNAPARTIALMETALAREA 8.956 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.346 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 17.334 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.809 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 15.576 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 54.656 LAYER METAL4 ;
  END iot_out[67]
  PIN iot_out[66] 
    ANTENNAPARTIALMETALAREA 8.454 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.589 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 7.94 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.93 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 12.87 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.185 LAYER METAL4 ;
  END iot_out[66]
  PIN iot_out[65] 
    ANTENNAPARTIALMETALAREA 9.53 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.355 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 6.866 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.171 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 9.21 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.375 LAYER METAL4 ;
  END iot_out[65]
  PIN iot_out[64] 
    ANTENNAPARTIALMETALAREA 9.12 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.92 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 15.974 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.049 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 13.044 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.794 LAYER METAL4 ;
  END iot_out[64]
  PIN iot_out[63] 
    ANTENNAPARTIALMETALAREA 8.792 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.772 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 15.208 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.368 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 19.594 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 68.719 LAYER METAL4 ;
  END iot_out[63]
  PIN iot_out[62] 
    ANTENNAPARTIALMETALAREA 9.848 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.468 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 10.628 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.338 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 19.574 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 68.649 LAYER METAL4 ;
  END iot_out[62]
  PIN iot_out[61] 
    ANTENNAPARTIALMETALAREA 11.006 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.521 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 9.974 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.049 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 18.168 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 63.728 LAYER METAL4 ;
  END iot_out[61]
  PIN iot_out[60] 
    ANTENNAPARTIALMETALAREA 7.224 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.284 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 11.64 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.88 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 26.092 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 91.462 LAYER METAL4 ;
  END iot_out[60]
  PIN iot_out[59] 
    ANTENNAPARTIALMETALAREA 6.896 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.136 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 14.4 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.54 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 26.43 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 92.645 LAYER METAL4 ;
  END iot_out[59]
  PIN iot_out[58] 
    ANTENNAPARTIALMETALAREA 8.372 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.302 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 15.924 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.874 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 25.21 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 88.375 LAYER METAL4 ;
  END iot_out[58]
  PIN iot_out[57] 
    ANTENNAPARTIALMETALAREA 9.602 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.607 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 14.472 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.792 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 24.092 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 84.462 LAYER METAL4 ;
  END iot_out[57]
  PIN iot_out[56] 
    ANTENNAPARTIALMETALAREA 7.47 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.145 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 11.272 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.592 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 21.694 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 76.069 LAYER METAL4 ;
  END iot_out[56]
  PIN iot_out[55] 
    ANTENNAPARTIALMETALAREA 6.568 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.988 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 15.32 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.76 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 23.13 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 81.095 LAYER METAL4 ;
  END iot_out[55]
  PIN iot_out[54] 
    ANTENNAPARTIALMETALAREA 8.874 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.059 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 14.686 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.541 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 20.906 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 73.311 LAYER METAL4 ;
  END iot_out[54]
  PIN iot_out[53] 
    ANTENNAPARTIALMETALAREA 9.12 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.92 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 11.364 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.914 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 24.472 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 85.792 LAYER METAL4 ;
  END iot_out[53]
  PIN iot_out[52] 
    ANTENNAPARTIALMETALAREA 8.208 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.728 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 14.492 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.862 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 20.168 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 70.728 LAYER METAL4 ;
  END iot_out[52]
  PIN iot_out[51] 
    ANTENNAPARTIALMETALAREA 7.224 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.284 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 11.732 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.202 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 23.776 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 83.356 LAYER METAL4 ;
  END iot_out[51]
  PIN iot_out[50] 
    ANTENNAPARTIALMETALAREA 6.814 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.849 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 12.458 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.743 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 25.918 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 90.853 LAYER METAL4 ;
  END iot_out[50]
  PIN iot_out[49] 
    ANTENNAPARTIALMETALAREA 6.978 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.423 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 10.996 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.626 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 27.998 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 98.133 LAYER METAL4 ;
  END iot_out[49]
  PIN iot_out[48] 
    ANTENNAPARTIALMETALAREA 9.274 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.459 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 11.19 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.305 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 26.05 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 91.315 LAYER METAL4 ;
  END iot_out[48]
  PIN iot_out[47] 
    ANTENNAPARTIALMETALAREA 7.798 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.293 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 8.614 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.289 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 26.328 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 92.288 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 1.162 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.207 LAYER METAL5 ;
  END iot_out[47]
  PIN iot_out[46] 
    ANTENNAPARTIALMETALAREA 9.038 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.633 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 7.766 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.321 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 31.832 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 111.552 LAYER METAL4 ;
  END iot_out[46]
  PIN iot_out[45] 
    ANTENNAPARTIALMETALAREA 9.11 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.885 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.45 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.715 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 28.512 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 99.932 LAYER METAL4 ;
  END iot_out[45]
  PIN iot_out[44] 
    ANTENNAPARTIALMETALAREA 10.012 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.042 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.266 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.071 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 31.596 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 110.726 LAYER METAL4 ;
  END iot_out[44]
  PIN iot_out[43] 
    ANTENNAPARTIALMETALAREA 9.11 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.885 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.15 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 32.19 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 112.805 LAYER METAL4 ;
  END iot_out[43]
  PIN iot_out[42] 
    ANTENNAPARTIALMETALAREA 7.306 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.571 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.898 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.783 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 32.468 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 113.778 LAYER METAL4 ;
  END iot_out[42]
  PIN iot_out[41] 
    ANTENNAPARTIALMETALAREA 8.792 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.772 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.646 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.901 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 32.94 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 115.43 LAYER METAL4 ;
  END iot_out[41]
  PIN iot_out[40] 
    ANTENNAPARTIALMETALAREA 15.526 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 54.341 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 8.206 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.861 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 27.844 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 97.594 LAYER METAL4 ;
  END iot_out[40]
  PIN iot_out[39] 
    ANTENNAPARTIALMETALAREA 8.454 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.589 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 13.286 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.641 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 35.562 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 124.607 LAYER METAL4 ;
  END iot_out[39]
  PIN iot_out[38] 
    ANTENNAPARTIALMETALAREA 7.634 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.719 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 13.03 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.745 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 35.254 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 123.529 LAYER METAL4 ;
  END iot_out[38]
  PIN iot_out[37] 
    ANTENNAPARTIALMETALAREA 5.994 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.979 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 13.204 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.354 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 36.742 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 128.737 LAYER METAL4 ;
  END iot_out[37]
  PIN iot_out[36] 
    ANTENNAPARTIALMETALAREA 7.47 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.145 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 22.926 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.381 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 34.322 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 120.267 LAYER METAL4 ;
  END iot_out[36]
  PIN iot_out[35] 
    ANTENNAPARTIALMETALAREA 24.374 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 85.309 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 41.364 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 144.914 LAYER METAL4 ;
  END iot_out[35]
  PIN iot_out[34] 
    ANTENNAPARTIALMETALAREA 21.132 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.962 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 40.564 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 142.114 LAYER METAL4 ;
  END iot_out[34]
  PIN iot_out[33] 
    ANTENNAPARTIALMETALAREA 19.292 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.522 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 31.288 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 109.648 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 7.674 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 26.999 LAYER METAL5 ;
  END iot_out[33]
  PIN iot_out[32] 
    ANTENNAPARTIALMETALAREA 26.076 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.266 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 38.064 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 133.364 LAYER METAL4 ;
  END iot_out[32]
  PIN iot_out[31] 
    ANTENNAPARTIALMETALAREA 28.708 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.478 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 33.892 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 118.762 LAYER METAL4 ;
  END iot_out[31]
  PIN iot_out[30] 
    ANTENNAPARTIALMETALAREA 31.642 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 110.747 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 32.776 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 114.856 LAYER METAL4 ;
  END iot_out[30]
  PIN iot_out[29] 
    ANTENNAPARTIALMETALAREA 30.14 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 105.49 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 31.874 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 111.699 LAYER METAL4 ;
  END iot_out[29]
  PIN iot_out[28] 
    ANTENNAPARTIALMETALAREA 8.058 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.203 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 15.914 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 55.839 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 23.794 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 83.419 LAYER METAL5 ;
  END iot_out[28]
  PIN iot_out[27] 
    ANTENNAPARTIALMETALAREA 9.08 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.78 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 31.626 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 110.831 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 24.53 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 85.995 LAYER METAL5 ;
  END iot_out[27]
  PIN iot_out[26] 
    ANTENNAPARTIALMETALAREA 9.54 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.39 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 12.306 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 43.211 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 25.633 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 89.8555 LAYER METAL5 ;
  END iot_out[26]
  PIN iot_out[25] 
    ANTENNAPARTIALMETALAREA 7.966 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.881 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 22.278 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 78.113 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 27.913 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 97.8355 LAYER METAL5 ;
  END iot_out[25]
  PIN iot_out[24] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.98 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 32.35 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 113.365 LAYER METAL5 ;
  END iot_out[24]
  PIN iot_out[23] 
    ANTENNAPARTIALMETALAREA 7.516 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.306 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 18.21 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 63.875 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 31.613 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 110.785 LAYER METAL5 ;
  END iot_out[23]
  PIN iot_out[22] 
    ANTENNAPARTIALMETALAREA 8.712 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.492 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 24.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 84.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 31.614 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 110.789 LAYER METAL5 ;
  END iot_out[22]
  PIN iot_out[21] 
    ANTENNAPARTIALMETALAREA 8.344 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.204 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 5.316 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.746 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 31.89 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 111.755 LAYER METAL5 ;
  END iot_out[21]
  PIN iot_out[20] 
    ANTENNAPARTIALMETALAREA 8.692 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.422 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.268 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 29.078 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 35.11 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 123.025 LAYER METAL5 ;
  END iot_out[20]
  PIN iot_out[19] 
    ANTENNAPARTIALMETALAREA 4.644 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.254 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.632 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.352 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 38.974 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 136.549 LAYER METAL5 ;
  END iot_out[19]
  PIN iot_out[18] 
    ANTENNAPARTIALMETALAREA 7.7 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.95 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 13.864 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 48.664 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 34.742 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 121.737 LAYER METAL5 ;
  END iot_out[18]
  PIN iot_out[17] 
    ANTENNAPARTIALMETALAREA 9.888 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.608 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 12.162 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 42.707 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 34.742 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 121.737 LAYER METAL5 ;
  END iot_out[17]
  PIN iot_out[16] 
    ANTENNAPARTIALMETALAREA 0.421 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4735 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.216 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 28.896 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 46.682 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 163.527 LAYER METAL5 ;
  END iot_out[16]
  PIN iot_out[15] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.98 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.55 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.065 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 47.05 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 164.815 LAYER METAL5 ;
  END iot_out[15]
  PIN iot_out[14] 
    ANTENNAPARTIALMETALAREA 8.16 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.56 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.491 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 34.282 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 120.127 LAYER METAL5 ;
  END iot_out[14]
  PIN iot_out[13] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.98 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.944 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.944 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 44.126 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 154.581 LAYER METAL5 ;
  END iot_out[13]
  PIN iot_out[12] 
    ANTENNAPARTIALMETALAREA 9.356 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.746 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 36.306 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 127.211 LAYER METAL5 ;
  END iot_out[12]
  PIN iot_out[11] 
    ANTENNAPARTIALMETALAREA 7.148 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.018 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.468 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.778 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 38.054 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 133.329 LAYER METAL5 ;
  END iot_out[11]
  PIN iot_out[10] 
    ANTENNAPARTIALMETALAREA 9.53 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.355 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 6.484 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.834 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 34.742 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 121.737 LAYER METAL5 ;
  END iot_out[10]
  PIN iot_out[9] 
    ANTENNAPARTIALMETALAREA 8.62 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.17 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.862 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.657 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 33.695 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 118.213 LAYER METAL5 ;
  END iot_out[9]
  PIN iot_out[8] 
    ANTENNAPARTIALMETALAREA 0.198 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.693 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.917 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 44.31 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 155.225 LAYER METAL5 ;
  END iot_out[8]
  PIN iot_out[7] 
    ANTENNAPARTIALMETALAREA 9.448 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.068 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.632 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.352 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 28.118 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 98.553 LAYER METAL5 ;
  END iot_out[7]
  PIN iot_out[6] 
    ANTENNAPARTIALMETALAREA 9.448 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.068 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.233 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 27.566 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 96.621 LAYER METAL5 ;
  END iot_out[6]
  PIN iot_out[5] 
    ANTENNAPARTIALMETALAREA 38.538 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 135.023 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 14.858 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 52.143 LAYER METAL4 ;
  END iot_out[5]
  PIN iot_out[4] 
    ANTENNAPARTIALMETALAREA 34.84 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 121.94 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 15.146 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 53.151 LAYER METAL4 ;
  END iot_out[4]
  PIN iot_out[3] 
    ANTENNAPARTIALMETALAREA 32.54 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 113.89 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 12.962 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.507 LAYER METAL4 ;
  END iot_out[3]
  PIN iot_out[2] 
    ANTENNAPARTIALMETALAREA 32.08 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 112.28 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 12.542 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 44.037 LAYER METAL4 ;
  END iot_out[2]
  PIN iot_out[1] 
    ANTENNAPARTIALMETALAREA 33.736 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 118.076 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 16.878 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 59.213 LAYER METAL4 ;
  END iot_out[1]
  PIN iot_out[0] 
    ANTENNAPARTIALMETALAREA 30.884 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 108.094 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.233 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 18.794 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 65.919 LAYER METAL4 ;
  END iot_out[0]
  PIN clk 
    ANTENNAPARTIALMETALAREA 0.09 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 21.034 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.759 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 46.224 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 161.924 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.3 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.33 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0754 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 17.2659 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 68.7692 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.91512 LAYER VIA56 ;
  END clk
  PIN rst 
    ANTENNAPARTIALMETALAREA 9.612 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.642 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 18.346 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.351 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 27.988 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 98.098 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 12.202 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 42.847 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8892 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 18.0893 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 62.9506 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.700321 LAYER VIA56 ;
  END rst
  PIN in_en 
    ANTENNAPARTIALMETALAREA 8.546 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.911 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 25.266 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 88.571 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 22.196 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 77.826 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6409 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 45.7724 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 161.963 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.21338 LAYER VIA45 ;
  END in_en
  PIN busy 
    ANTENNAPARTIALMETALAREA 8.618 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.163 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 10.351 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.3685 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3646 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 22.884 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 80.234 LAYER METAL4 ;
  END busy
  PIN valid 
    ANTENNAPARTIALMETALAREA 7.716 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.006 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 9.248 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.508 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 27.968 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 98.028 LAYER METAL4 ;
  END valid
END IOTDF

END LIBRARY
