

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO IOTDF 
  PIN clk 
    ANTENNAPARTIALMETALAREA 0.09 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.61 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.275 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 23.018 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 80.703 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 381.452 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1339.12 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.02849 LAYER VIA45 ;
  END clk
  PIN rst 
    ANTENNAPARTIALMETALAREA 8.984 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.584 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8268 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 11.0766 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 38.9204 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.0436623 LAYER VIA23 ;
  END rst
  PIN in_en 
    ANTENNAPARTIALMETALAREA 7.204 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.214 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 31.338 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 109.823 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 23.14 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 81.13 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4927 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 58.3613 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 204.67 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.381872 LAYER VIA45 ;
  END in_en
  PIN iot_in[7] 
    ANTENNAPARTIALMETALAREA 18.541 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 64.8935 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 6.816 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.996 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 68.0233 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 240.788 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.68566 LAYER VIA34 ;
  END iot_in[7]
  PIN iot_in[6] 
    ANTENNAPARTIALMETALAREA 16.03 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 56.105 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 8.554 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.079 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 101.623 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 358.386 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.68566 LAYER VIA34 ;
  END iot_in[6]
  PIN iot_in[5] 
    ANTENNAPARTIALMETALAREA 0.072 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.252 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.054 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.969 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.584 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.684 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 82.8381 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 293.97 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.02849 LAYER VIA45 ;
  END iot_in[5]
  PIN iot_in[4] 
    ANTENNAPARTIALMETALAREA 7.636 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.726 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.794 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.919 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.36 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 29.4 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 90.2455 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 319.896 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.02849 LAYER VIA45 ;
  END iot_in[4]
  PIN iot_in[3] 
    ANTENNAPARTIALMETALAREA 12.932 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 45.542 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 124.737 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 439.288 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.34283 LAYER VIA23 ;
  END iot_in[3]
  PIN iot_in[2] 
    ANTENNAPARTIALMETALAREA 12.481 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 43.9635 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 120.454 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 424.297 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.34283 LAYER VIA23 ;
  END iot_in[2]
  PIN iot_in[1] 
    ANTENNAPARTIALMETALAREA 9.943 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.0805 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 96.3519 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 339.938 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.34283 LAYER VIA23 ;
  END iot_in[1]
  PIN iot_in[0] 
    ANTENNAPARTIALMETALAREA 12.565 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 44.2575 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 121.252 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 427.089 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.34283 LAYER VIA23 ;
  END iot_in[0]
  PIN fn_sel[2] 
    ANTENNAPARTIALMETALAREA 9.916 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.706 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.83 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.545 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 26.9831 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 95.8188 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 4.404 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.554 LAYER METAL4 ;
    ANTENNAGATEAREA 0.3952 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 38.1268 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 135.176 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.04508 LAYER VIA45 ;
  END fn_sel[2]
  PIN fn_sel[1] 
    ANTENNAPARTIALMETALAREA 6.997 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.4895 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.082 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.427 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 4.404 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.554 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4121 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 21.1471 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 75.051 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.73558 LAYER VIA45 ;
  END fn_sel[1]
  PIN fn_sel[0] 
    ANTENNAPARTIALMETALAREA 9.826 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.391 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.622 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.817 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2561 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 7.45041 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 26.802 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.422882 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.03 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.745 LAYER METAL4 ;
    ANTENNAGATEAREA 1.3533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 12.6215 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 44.7979 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.649996 LAYER VIA45 ;
  END fn_sel[0]
  PIN busy 
    ANTENNADIFFAREA 0.3646 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 9.999 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.1365 LAYER METAL2 ;
  END busy
  PIN valid 
    ANTENNAPARTIALMETALAREA 0.089 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3115 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 4.474 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.799 LAYER METAL3 ;
  END valid
  PIN iot_out[127] 
    ANTENNAPARTIALMETALAREA 6.295 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.0325 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.99 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.105 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 7.028 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 24.738 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 22.2408 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 79.4772 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[127]
  PIN iot_out[126] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 13.863 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 48.8005 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 30.111 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 104.824 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.322898 LAYER VIA23 ;
  END iot_out[126]
  PIN iot_out[125] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 13.473 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 47.2955 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 27.1566 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 94.537 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[125]
  PIN iot_out[124] 
    ANTENNAPARTIALMETALAREA 8.662 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.317 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.338 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.323 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 16.7827 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 58.1731 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.395214 LAYER VIA34 ;
  END iot_out[124]
  PIN iot_out[123] 
    ANTENNAPARTIALMETALAREA 8.189 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.6615 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.416 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.736 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 18.5887 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 65.1672 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.455233 LAYER VIA34 ;
  END iot_out[123]
  PIN iot_out[122] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 12.241 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 42.9835 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 26.1735 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 90.8722 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.322898 LAYER VIA23 ;
  END iot_out[122]
  PIN iot_out[121] 
    ANTENNAPARTIALMETALAREA 10.664 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 37.464 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 28.3025 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 98.8352 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.319568 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.518 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.953 LAYER METAL3 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 29.2512 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 102.412 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[121]
  PIN iot_out[120] 
    ANTENNAPARTIALMETALAREA 9.595 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.7225 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.234 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 41.7171 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 145.98 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.308547 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.794 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.919 LAYER METAL3 ;
    ANTENNAGATEAREA 0.234 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 45.1103 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 158.454 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.462821 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.026 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.231 LAYER METAL4 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 49.1688 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 172.939 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.968694 LAYER VIA45 ;
  END iot_out[120]
  PIN iot_out[119] 
    ANTENNAPARTIALMETALAREA 8.929 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.3915 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.234 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 39.5192 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 138.196 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.308547 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.692 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.702 LAYER METAL3 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 44.4496 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 155.965 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.466743 LAYER VIA34 ;
  END iot_out[119]
  PIN iot_out[118] 
    ANTENNAPARTIALMETALAREA 9.614 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.789 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.234 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 51.8158 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 178.731 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.462821 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.794 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.919 LAYER METAL3 ;
    ANTENNAGATEAREA 0.3458 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 54.1119 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 187.172 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.750192 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.748 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.258 LAYER METAL4 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 61.6199 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 213.731 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.750192 LAYER VIA45 ;
  END iot_out[118]
  PIN iot_out[117] 
    ANTENNAPARTIALMETALAREA 6.162 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.567 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.542 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.037 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 8.708 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 30.618 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 26.8176 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 94.3073 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.367567 LAYER VIA45 ;
  END iot_out[117]
  PIN iot_out[116] 
    ANTENNAPARTIALMETALAREA 7.662 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.817 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.29 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.155 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 10.256 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.036 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 34.9136 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 121.506 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.467529 LAYER VIA45 ;
  END iot_out[116]
  PIN iot_out[115] 
    ANTENNAPARTIALMETALAREA 7.924 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.734 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 11.19 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.305 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 11.004 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.654 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 32.7501 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 115.003 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.433684 LAYER VIA45 ;
  END iot_out[115]
  PIN iot_out[114] 
    ANTENNAPARTIALMETALAREA 6.659 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.3065 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 13.674 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.999 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 16.526 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 58.121 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 40.6671 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 142.487 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[114]
  PIN iot_out[113] 
    ANTENNAPARTIALMETALAREA 6.057 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.1995 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 17.794 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.419 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 18.987 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 66.5945 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 38.9677 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 138.021 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[113]
  PIN iot_out[112] 
    ANTENNAPARTIALMETALAREA 6.447 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.5645 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 20.85 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.115 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 14.332 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 50.442 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 34.8751 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 122.661 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.612161 LAYER VIA45 ;
  END iot_out[112]
  PIN iot_out[111] 
    ANTENNAPARTIALMETALAREA 7.236 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.326 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 23.334 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 81.809 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 13.594 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 47.859 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 51.9851 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 183.439 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.838232 LAYER VIA45 ;
  END iot_out[111]
  PIN iot_out[110] 
    ANTENNAPARTIALMETALAREA 8.074 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.259 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 27.72 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 97.16 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 17.284 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 60.774 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 45.143 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 158.151 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.603653 LAYER VIA45 ;
  END iot_out[110]
  PIN iot_out[109] 
    ANTENNAPARTIALMETALAREA 7.594 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.579 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 31.594 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 110.719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 16.468 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 57.778 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 38.0657 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 134.544 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[109]
  PIN iot_out[108] 
    ANTENNAPARTIALMETALAREA 6.814 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.849 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 37.042 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 129.787 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 12.932 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.402 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 46.6742 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 164.597 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.542981 LAYER VIA45 ;
  END iot_out[108]
  PIN iot_out[107] 
    ANTENNAPARTIALMETALAREA 23.064 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.724 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 43.762 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 153.307 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 88.9935 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 311.923 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.433684 LAYER VIA45 ;
  END iot_out[107]
  PIN iot_out[106] 
    ANTENNAPARTIALMETALAREA 21.405 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.9175 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 38.864 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 136.164 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 92.517 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 324.796 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.778313 LAYER VIA45 ;
  END iot_out[106]
  PIN iot_out[105] 
    ANTENNAPARTIALMETALAREA 21.586 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 75.551 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 34.262 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 120.057 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 74.2374 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 260.896 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.536782 LAYER VIA45 ;
  END iot_out[105]
  PIN iot_out[104] 
    ANTENNAPARTIALMETALAREA 18.823 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.8805 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 31.924 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 111.874 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 81.8499 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 286.569 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.371221 LAYER VIA45 ;
  END iot_out[104]
  PIN iot_out[103] 
    ANTENNAPARTIALMETALAREA 20.016 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 70.056 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 28.388 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 99.498 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 70.6837 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 247.963 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.528938 LAYER VIA45 ;
  END iot_out[103]
  PIN iot_out[102] 
    ANTENNAPARTIALMETALAREA 20.923 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.2305 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 24.042 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 84.287 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 66.2496 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 232.318 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.718112 LAYER VIA45 ;
  END iot_out[102]
  PIN iot_out[101] 
    ANTENNAPARTIALMETALAREA 25.64 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.74 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 20.978 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 73.563 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 48.6264 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 171.171 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.536782 LAYER VIA45 ;
  END iot_out[101]
  PIN iot_out[100] 
    ANTENNAPARTIALMETALAREA 23.432 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 82.012 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 19.92 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 69.86 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 55.3201 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 195.49 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.968694 LAYER VIA45 ;
  END iot_out[100]
  PIN iot_out[99] 
    ANTENNAPARTIALMETALAREA 18.214 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.749 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 13.178 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 46.263 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 4.464 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.764 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 24.2589 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 84.9963 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.598977 LAYER VIA56 ;
  END iot_out[99]
  PIN iot_out[98] 
    ANTENNAPARTIALMETALAREA 11.704 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.964 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 10.638 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 37.373 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 56.1272 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 196.763 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.539845 LAYER VIA56 ;
  END iot_out[98]
  PIN iot_out[97] 
    ANTENNAPARTIALMETALAREA 0.254 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.889 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.632 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.352 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 22.506 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 78.911 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 53.9367 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 189.224 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.433684 LAYER VIA56 ;
  END iot_out[97]
  PIN iot_out[96] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.714 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.639 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 21.218 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 74.403 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 56.5206 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 197.98 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.676321 LAYER VIA56 ;
  END iot_out[96]
  PIN iot_out[95] 
    ANTENNAPARTIALMETALAREA 18.832 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.912 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.584 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.684 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 20.7403 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 73.5692 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.536782 LAYER VIA45 ;
  END iot_out[95]
  PIN iot_out[94] 
    ANTENNADIFFAREA 0.4012 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.928 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.248 LAYER METAL3 ;
  END iot_out[94]
  PIN iot_out[93] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.13 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.595 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 27.7302 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 97.7845 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.645796 LAYER VIA34 ;
  END iot_out[93]
  PIN iot_out[92] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 4.598 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.233 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 39.2405 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 131.627 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.617094 LAYER VIA34 ;
  END iot_out[92]
  PIN iot_out[91] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.55 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.925 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 26.4012 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 92.0461 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.455233 LAYER VIA34 ;
  END iot_out[91]
  PIN iot_out[90] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.721 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.5235 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 27.2526 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 95.5227 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[90]
  PIN iot_out[89] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.248 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.008 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 29.2976 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 102.677 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[89]
  PIN iot_out[88] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 6.306 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.211 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 44.3867 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 148.971 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.492449 LAYER VIA34 ;
  END iot_out[88]
  PIN iot_out[87] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.668 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.118 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 45.6234 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 159.572 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.910467 LAYER VIA34 ;
  END iot_out[87]
  PIN iot_out[86] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 11.568 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.628 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 28.4487 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 99.7075 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.367567 LAYER VIA34 ;
  END iot_out[86]
  PIN iot_out[85] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.572 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.142 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 34.0703 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 119.905 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.547184 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 0.796 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.926 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 35.5282 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 125.264 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[85]
  PIN iot_out[84] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.644 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 32.8451 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 115.359 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[84]
  PIN iot_out[83] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.638 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.373 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 30.9096 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 109.117 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[83]
  PIN iot_out[82] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.94 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.71 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 28.1501 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 99.4389 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[82]
  PIN iot_out[81] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 11.782 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.377 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.312 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 39.8107 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 140.089 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.58637 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 0.878 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.213 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 41.4188 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 145.974 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.58637 LAYER VIA45 ;
  END iot_out[81]
  PIN iot_out[80] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 11.599 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.7365 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 24.327 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 85.1775 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[80]
  PIN iot_out[79] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 11.368 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.928 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 28.4729 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 99.4796 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.351038 LAYER VIA34 ;
  END iot_out[79]
  PIN iot_out[78] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.311 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.7285 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 29.4752 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 103.446 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[78]
  PIN iot_out[77] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.957 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.4895 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 25.7027 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 90.7681 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.455233 LAYER VIA34 ;
  END iot_out[77]
  PIN iot_out[76] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.376 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.096 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 80.0518 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 280.997 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[76]
  PIN iot_out[75] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 15.651 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.9185 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 40.0441 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 138.653 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.351038 LAYER VIA34 ;
  END iot_out[75]
  PIN iot_out[74] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 14.796 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.926 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 50.368 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 176.205 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.455233 LAYER VIA34 ;
  END iot_out[74]
  PIN iot_out[73] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 17.167 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.3645 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 35.1525 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 123.691 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[73]
  PIN iot_out[72] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.002 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.647 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 116.567 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 408.545 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.68285 LAYER VIA34 ;
  END iot_out[72]
  PIN iot_out[71] 
    ANTENNAPARTIALMETALAREA 24.864 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 87.024 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 11.178 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.263 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 33.6391 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 118.368 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[71]
  PIN iot_out[70] 
    ANTENNAPARTIALMETALAREA 21.113 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 73.8955 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 6.58 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.17 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.358 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.893 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 11.3708 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 41.6439 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[70]
  PIN iot_out[69] 
    ANTENNAPARTIALMETALAREA 21.039 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 73.7765 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 6.499 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.8865 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 21.3762 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 75.5386 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[69]
  PIN iot_out[68] 
    ANTENNAPARTIALMETALAREA 19.935 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 69.7725 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 5.926 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.881 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 12.9014 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 45.714 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[68]
  PIN iot_out[67] 
    ANTENNAPARTIALMETALAREA 16.358 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 57.253 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.234 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 72.2038 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 251.76 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.308547 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 3.888 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.888 LAYER METAL3 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 79.3247 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 277.196 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.466743 LAYER VIA34 ;
  END iot_out[67]
  PIN iot_out[66] 
    ANTENNAPARTIALMETALAREA 16.825 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.8875 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.234 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 72.5615 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 253.512 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.308547 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.266 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.071 LAYER METAL3 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 76.7117 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 268.294 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.417155 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 1.534 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.509 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 79.5212 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 278.383 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.417155 LAYER VIA45 ;
  END iot_out[66]
  PIN iot_out[65] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 16.295 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 57.0325 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 32.2041 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 111.66 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[65]
  PIN iot_out[64] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 15.762 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 55.167 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.89 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.255 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 8.54474 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 29.8393 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.30145 LAYER VIA34 ;
  END iot_out[64]
  PIN iot_out[63] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 13.436 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 47.306 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3874 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 51.6515 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 176.976 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.56385 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.426 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.631 LAYER METAL3 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 52.4318 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 179.963 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.56385 LAYER VIA34 ;
  END iot_out[63]
  PIN iot_out[62] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 14.968 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 52.668 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 32.4142 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 112.428 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA23 ;
  END iot_out[62]
  PIN iot_out[61] 
    ANTENNAPARTIALMETALAREA 12.832 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 45.052 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 36.248 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 123.468 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.374664 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.977 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5595 LAYER METAL3 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 38.0374 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 129.988 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.374664 LAYER VIA34 ;
  END iot_out[61]
  PIN iot_out[60] 
    ANTENNAPARTIALMETALAREA 10.127 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.4445 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.37 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.935 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 9.27473 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 32.7909 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.417155 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.272 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.092 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 13.4359 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 47.6114 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.417155 LAYER VIA45 ;
  END iot_out[60]
  PIN iot_out[59] 
    ANTENNAPARTIALMETALAREA 7.97 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.895 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 3.762 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.587 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 18.976 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 66.9855 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.466743 LAYER VIA34 ;
  END iot_out[59]
  PIN iot_out[58] 
    ANTENNAPARTIALMETALAREA 10.308 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.078 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.714 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.139 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 13.0977 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 45.8168 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.30145 LAYER VIA34 ;
  END iot_out[58]
  PIN iot_out[57] 
    ANTENNAPARTIALMETALAREA 12.63 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 44.345 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 32.1037 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 109.907 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.374664 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.978 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.563 LAYER METAL3 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 33.8949 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 116.432 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.374664 LAYER VIA34 ;
  END iot_out[57]
  PIN iot_out[56] 
    ANTENNAPARTIALMETALAREA 8.466 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.631 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.502 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.037 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 11.6774 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 41.3607 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.50347 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.174 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.249 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 18.3383 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 65.1449 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[56]
  PIN iot_out[55] 
    ANTENNAPARTIALMETALAREA 9.236 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.326 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.334 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.309 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 11.414 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 40.089 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 30.3773 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 106.97 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.433684 LAYER VIA45 ;
  END iot_out[55]
  PIN iot_out[54] 
    ANTENNAPARTIALMETALAREA 7.486 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.201 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.886 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.241 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 12.87 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.185 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 39.7302 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 140.377 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.748967 LAYER VIA45 ;
  END iot_out[54]
  PIN iot_out[53] 
    ANTENNAPARTIALMETALAREA 0.085 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2975 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.358 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 22.852 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 80.122 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 67.9239 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 239.368 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[53]
  PIN iot_out[52] 
    ANTENNAPARTIALMETALAREA 0.313 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0955 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.334 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.309 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 23.546 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 82.691 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 66.118 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 233.304 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[52]
  PIN iot_out[51] 
    ANTENNAPARTIALMETALAREA 8.466 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.631 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.358 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 11.968 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 42.028 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 41.0298 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 144.399 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.536782 LAYER VIA45 ;
  END iot_out[51]
  PIN iot_out[50] 
    ANTENNAPARTIALMETALAREA 7.624 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.684 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.738 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.223 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 17.318 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 60.753 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 39.9373 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 141.626 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[50]
  PIN iot_out[49] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2135 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.542 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.037 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 23.878 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 83.713 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 49.2956 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 173.173 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.521351 LAYER VIA45 ;
  END iot_out[49]
  PIN iot_out[48] 
    ANTENNAPARTIALMETALAREA 0.093 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3255 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.254 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.529 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 20.638 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 72.373 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 50.5939 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 177.992 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.536782 LAYER VIA45 ;
  END iot_out[48]
  PIN iot_out[47] 
    ANTENNAPARTIALMETALAREA 8.837 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.0695 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.886 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.241 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 7.37788 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 25.9557 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.411519 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.42 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.11 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 19.3338 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 69.1026 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[47]
  PIN iot_out[46] 
    ANTENNAPARTIALMETALAREA 8.162 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.567 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 11.65 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.915 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 34.3269 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 120.527 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.411519 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 5.162 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.207 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 43.7811 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 153.873 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[46]
  PIN iot_out[45] 
    ANTENNAPARTIALMETALAREA 10.455 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.7325 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.234 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 45.3393 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 158.832 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.308547 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.794 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.919 LAYER METAL3 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 47.3617 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 166.267 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.547184 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.338 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.823 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 53.4753 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 187.921 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[45]
  PIN iot_out[44] 
    ANTENNAPARTIALMETALAREA 7.37 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.795 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 14.554 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.219 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.234 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 70.4632 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 247.962 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.617094 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 1.39 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.005 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 73.009 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 257.129 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.617094 LAYER VIA45 ;
  END iot_out[44]
  PIN iot_out[43] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 14.201 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.8435 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 27.0861 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 94.6819 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[43]
  PIN iot_out[42] 
    ANTENNAPARTIALMETALAREA 7.729 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.0515 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.732 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.342 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 31.5026 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 110.448 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.367567 LAYER VIA34 ;
  END iot_out[42]
  PIN iot_out[41] 
    ANTENNAPARTIALMETALAREA 9.712 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.132 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 25.8016 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 90.3318 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.319568 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL3 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 26.1684 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 91.9721 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.411519 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 4.486 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.841 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 34.3845 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 120.985 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[41]
  PIN iot_out[40] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 14.162 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.847 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 30.9788 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 107.363 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA23 ;
  END iot_out[40]
  PIN iot_out[39] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 14.644 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 51.534 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 30.8925 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 107.334 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA23 ;
  END iot_out[39]
  PIN iot_out[38] 
    ANTENNAPARTIALMETALAREA 9.689 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.0515 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 25.7431 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 90.1268 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.319568 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.15 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER METAL3 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 26.1251 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 91.8206 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.411519 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.092 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 31.7881 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 111.898 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[38]
  PIN iot_out[37] 
    ANTENNAPARTIALMETALAREA 9.151 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.0285 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 13.562 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.607 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 36.5674 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 127.98 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.411519 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.928 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.388 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 41.9301 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 147.005 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[37]
  PIN iot_out[36] 
    ANTENNAPARTIALMETALAREA 9.433 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.1555 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 25.1009 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 87.8445 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.319568 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.987 LAYER METAL3 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 25.7173 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 90.3585 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.411519 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.272 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.092 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 29.8785 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 105.179 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[36]
  PIN iot_out[35] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.542 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.037 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 31.57 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 110.26 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.293734 LAYER VIA34 ;
  END iot_out[35]
  PIN iot_out[34] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.785 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.8875 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 44.3854 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 155.282 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.367567 LAYER VIA34 ;
  END iot_out[34]
  PIN iot_out[33] 
    ANTENNAPARTIALMETALAREA 10.41 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.575 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 44.3039 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 155.446 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.50347 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.42 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.11 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 50.5677 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 177.626 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[33]
  PIN iot_out[32] 
    ANTENNAPARTIALMETALAREA 8.319 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.2565 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 37.7375 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 132.82 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.50347 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.928 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.388 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 43.1001 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 151.846 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[32]
  PIN iot_out[31] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.892 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.262 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 24.4833 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 85.4064 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.30145 LAYER VIA34 ;
  END iot_out[31]
  PIN iot_out[30] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.739 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.7265 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 1.206 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.361 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 7.19953 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 25.637 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.367567 LAYER VIA45 ;
  END iot_out[30]
  PIN iot_out[29] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 9.924 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.014 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.682 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.527 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 10.3431 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 36.4902 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.536782 LAYER VIA45 ;
  END iot_out[29]
  PIN iot_out[28] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 10.856 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.136 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 38.9779 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 136.548 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.351038 LAYER VIA34 ;
  END iot_out[28]
  PIN iot_out[27] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 14.262 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.337 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 56.0547 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 197.564 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.774801 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.19 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.805 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 60.0657 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 211.859 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.774801 LAYER VIA45 ;
  END iot_out[27]
  PIN iot_out[26] 
    ANTENNAPARTIALMETALAREA 0.174 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.609 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 13.858 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 48.643 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 48.6379 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 171.724 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.602899 LAYER VIA56 ;
  END iot_out[26]
  PIN iot_out[25] 
    ANTENNAPARTIALMETALAREA 15.404 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.914 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 7.356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 25.886 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 19.9622 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 70.8459 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.536782 LAYER VIA45 ;
  END iot_out[25]
  PIN iot_out[24] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 17.55 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.565 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.256 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.536 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 13.6454 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 48.9485 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.536782 LAYER VIA45 ;
  END iot_out[24]
  PIN iot_out[23] 
    ANTENNAPARTIALMETALAREA 9.11 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.885 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.714 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.639 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 9.994 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 35.119 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 41.392 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 146.45 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.815084 LAYER VIA56 ;
  END iot_out[23]
  PIN iot_out[22] 
    ANTENNAPARTIALMETALAREA 0.248 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.868 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.19 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.805 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 17.446 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 61.201 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 44.3857 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 155.756 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.602899 LAYER VIA56 ;
  END iot_out[22]
  PIN iot_out[21] 
    ANTENNAPARTIALMETALAREA 4.596 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.086 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 14.778 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 51.863 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 40.648 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 142.839 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.602899 LAYER VIA56 ;
  END iot_out[21]
  PIN iot_out[20] 
    ANTENNAPARTIALMETALAREA 8.675 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.3625 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.108 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.518 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 12.55 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 44.065 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 33.2018 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 118.753 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.94133 LAYER VIA56 ;
  END iot_out[20]
  PIN iot_out[19] 
    ANTENNAPARTIALMETALAREA 0.236 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.826 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 18.09 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 63.455 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 48.1145 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 169.315 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.602899 LAYER VIA56 ;
  END iot_out[19]
  PIN iot_out[18] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 22.196 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 77.826 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 48.879 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 171.636 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.68285 LAYER VIA34 ;
  END iot_out[18]
  PIN iot_out[17] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 21.88 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.86 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 45.6329 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 160.905 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[17]
  PIN iot_out[16] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 21.628 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 75.698 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 45.1694 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 158.232 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[16]
  PIN iot_out[15] 
    ANTENNAPARTIALMETALAREA 9.106 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.011 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.584 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.684 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 18.5995 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 66.0139 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[15]
  PIN iot_out[14] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 10.522 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.107 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 48.1325 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 169.675 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.94133 LAYER VIA34 ;
  END iot_out[14]
  PIN iot_out[13] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.376 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.456 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 25.2064 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 88.7814 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[13]
  PIN iot_out[12] 
    ANTENNAPARTIALMETALAREA 10.99 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.745 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 25.9835 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 91.9205 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.772115 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 1.452 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.222 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 28.6428 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 101.485 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.772115 LAYER VIA45 ;
  END iot_out[12]
  PIN iot_out[11] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.784 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 27.3884 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 96.1486 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[11]
  PIN iot_out[10] 
    ANTENNAPARTIALMETALAREA 10.826 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.171 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 27.4364 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 96.6846 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.536782 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 0.96 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 29.1946 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 103.095 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.536782 LAYER VIA45 ;
  END iot_out[10]
  PIN iot_out[9] 
    ANTENNAPARTIALMETALAREA 10.198 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.833 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3926 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 29.4733 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 104.065 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.547184 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 1.452 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.222 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 32.1327 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 113.63 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[9]
  PIN iot_out[8] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.628 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.118 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 30.1827 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 106.874 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[8]
  PIN iot_out[7] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 11.64 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.02 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 28.0021 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 98.0573 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.367567 LAYER VIA34 ;
  END iot_out[7]
  PIN iot_out[6] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.112 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.032 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 28.1424 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 99.2203 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[6]
  PIN iot_out[5] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.321 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.9035 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 33.1911 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 116.947 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[5]
  PIN iot_out[4] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.989 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.2415 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 29.7117 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 104.838 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[4]
  PIN iot_out[3] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 11.075 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.1825 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 66.2788 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 233.048 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[3]
  PIN iot_out[2] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 11.318 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.893 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 26.7664 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 94.214 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[2]
  PIN iot_out[1] 
    ANTENNAPARTIALMETALAREA 11.143 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.1405 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 120.066 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 421.611 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.94133 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.986 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.731 LAYER METAL4 ;
    ANTENNAGATEAREA 0.546 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 125.535 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 441.265 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.94133 LAYER VIA45 ;
  END iot_out[1]
  PIN iot_out[0] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.248 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.508 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 122.6 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 429.827 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.968694 LAYER VIA34 ;
  END iot_out[0]
END IOTDF

END LIBRARY
