

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO IOTDF 
  PIN iot_in[7] 
    ANTENNAPARTIALMETALAREA 13.301 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 46.5535 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 8.748 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.758 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 87.8903 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 310.323 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.68566 LAYER VIA34 ;
  END iot_in[7]
  PIN iot_in[6] 
    ANTENNAPARTIALMETALAREA 5.91 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.685 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.842 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.087 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.872 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 31.192 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 112.544 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 397.939 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.02849 LAYER VIA45 ;
  END iot_in[6]
  PIN iot_in[5] 
    ANTENNAPARTIALMETALAREA 0.086 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.301 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.987 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 10.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 35.644 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 126.39 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 446.401 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.02849 LAYER VIA45 ;
  END iot_in[5]
  PIN iot_in[4] 
    ANTENNAPARTIALMETALAREA 0.083 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2905 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.278 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.613 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.852 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 31.122 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 90.5304 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 320.893 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.02849 LAYER VIA45 ;
  END iot_in[4]
  PIN iot_in[3] 
    ANTENNAPARTIALMETALAREA 7.786 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.391 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 75.8675 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 266.914 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.34283 LAYER VIA23 ;
  END iot_in[3]
  PIN iot_in[2] 
    ANTENNAPARTIALMETALAREA 11.391 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 40.0085 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 110.103 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 386.738 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.34283 LAYER VIA23 ;
  END iot_in[2]
  PIN iot_in[1] 
    ANTENNAPARTIALMETALAREA 0.074 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.259 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.987 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 12.85 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.115 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 128.213 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 452.783 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.02849 LAYER VIA45 ;
  END iot_in[1]
  PIN iot_in[0] 
    ANTENNAPARTIALMETALAREA 0.071 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2485 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.987 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 13.772 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 48.342 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 139.049 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 490.708 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.02849 LAYER VIA45 ;
  END iot_in[0]
  PIN fn_sel[2] 
    ANTENNAPARTIALMETALAREA 8.196 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.686 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.154 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1586 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 16.0451 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 57.5927 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.68285 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.494 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.009 LAYER METAL4 ;
    ANTENNAGATEAREA 1.1206 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 30.9149 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 111.128 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.08553 LAYER VIA45 ;
  END fn_sel[2]
  PIN fn_sel[1] 
    ANTENNAPARTIALMETALAREA 8.511 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.7885 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 51.4332 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 174.456 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.741874 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.702 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.597 LAYER METAL3 ;
    ANTENNAGATEAREA 0.3744 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 53.3082 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 181.393 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.741874 LAYER VIA34 ;
  END fn_sel[1]
  PIN fn_sel[0] 
    ANTENNAPARTIALMETALAREA 9.245 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.4975 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2158 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 45.9916 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 158.841 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.74581 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.518 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.953 LAYER METAL3 ;
    ANTENNAGATEAREA 0.4719 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 47.0893 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 162.979 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.74581 LAYER VIA34 ;
  END fn_sel[0]
  PIN iot_out[127] 
    ANTENNAPARTIALMETALAREA 6.043 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.1505 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 3.256 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.536 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 29.941 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 106.884 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[127]
  PIN iot_out[126] 
    ANTENNAPARTIALMETALAREA 7.679 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.8765 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.22 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.55 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 26.0443 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 93.4459 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[126]
  PIN iot_out[125] 
    ANTENNAPARTIALMETALAREA 0.148 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.518 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.953 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 9.16 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.2 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 66.7005 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 235.954 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[125]
  PIN iot_out[124] 
    ANTENNAPARTIALMETALAREA 0.15 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 9.672 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.992 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 75.8879 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 267.898 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[124]
  PIN iot_out[123] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 7.098 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.983 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 47.3481 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 166.184 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[123]
  PIN iot_out[122] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 7.09 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.955 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 47.296 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 166.001 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[122]
  PIN iot_out[121] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 7.092 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.962 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 47.309 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 166.047 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[121]
  PIN iot_out[120] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 7.643 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.0305 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 50.7291 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 179.141 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[120]
  PIN iot_out[119] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 7.646 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.761 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.61 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.275 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 9.00163 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 33.0952 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[119]
  PIN iot_out[118] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 8.237 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.8295 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 58.0962 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 202.089 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[118]
  PIN iot_out[117] 
    ANTENNAPARTIALMETALAREA 0.074 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.259 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.806 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.461 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 9.672 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.992 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 74.0887 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 261.601 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[117]
  PIN iot_out[116] 
    ANTENNAPARTIALMETALAREA 3.941 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.7935 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.91 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.325 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 8.596 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 30.226 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 75.1033 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 265.364 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[116]
  PIN iot_out[115] 
    ANTENNAPARTIALMETALAREA 4.354 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.239 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.106 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.511 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 10.984 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.584 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 93.263 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 328.391 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[115]
  PIN iot_out[114] 
    ANTENNAPARTIALMETALAREA 7.626 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.691 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 6.846 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.101 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 9.406 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.061 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 78.7063 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 277.436 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[114]
  PIN iot_out[113] 
    ANTENNAPARTIALMETALAREA 6.809 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.8315 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 15.116 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.046 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 9.426 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.131 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 75.8393 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 267.638 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[113]
  PIN iot_out[112] 
    ANTENNAPARTIALMETALAREA 6.331 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.1585 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 15.474 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.299 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 11.968 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 42.028 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 94.6268 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 332.95 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[112]
  PIN iot_out[111] 
    ANTENNAPARTIALMETALAREA 4.602 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.107 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 16.526 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.981 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 13.556 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 47.586 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 107.778 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 380.428 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[111]
  PIN iot_out[110] 
    ANTENNAPARTIALMETALAREA 4.933 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2655 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 21.218 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.403 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 13.926 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 48.881 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 100.541 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 353.983 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[110]
  PIN iot_out[109] 
    ANTENNAPARTIALMETALAREA 5.92 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.72 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 23.058 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.843 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 13.69 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 48.055 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 107.933 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 379.857 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[109]
  PIN iot_out[108] 
    ANTENNAPARTIALMETALAREA 5.338 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.683 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 28.578 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.163 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 12.614 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 44.289 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 103.393 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 363.841 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[108]
  PIN iot_out[107] 
    ANTENNAPARTIALMETALAREA 19.568 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 68.488 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 29.608 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 103.768 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 206.395 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 724.355 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[107]
  PIN iot_out[106] 
    ANTENNAPARTIALMETALAREA 20.479 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.6765 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 26.954 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 94.479 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 181.846 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 638.752 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[106]
  PIN iot_out[105] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 20.395 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.5225 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 138.539 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 486.066 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[105]
  PIN iot_out[104] 
    ANTENNAPARTIALMETALAREA 18.718 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.513 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 20.66 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 72.45 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 148.676 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 522.867 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[104]
  PIN iot_out[103] 
    ANTENNAPARTIALMETALAREA 18.067 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.2345 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 18.24 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 63.98 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 140.462 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 494.119 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[103]
  PIN iot_out[102] 
    ANTENNAPARTIALMETALAREA 21.686 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 75.901 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 10.246 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.001 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 76.7744 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 271.001 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[102]
  PIN iot_out[101] 
    ANTENNAPARTIALMETALAREA 16.465 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.6275 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 8.278 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 29.113 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 97.322 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 342.918 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[101]
  PIN iot_out[100] 
    ANTENNAPARTIALMETALAREA 13.546 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.411 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 5.684 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.034 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 84.3015 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 297.557 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[100]
  PIN iot_out[99] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 18.887 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.2445 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 0.386 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.491 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 5.50978 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 21.575 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[99]
  PIN iot_out[98] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 16.116 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.406 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 132.029 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 462.566 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[98]
  PIN iot_out[97] 
    ANTENNAPARTIALMETALAREA 9.807 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.3245 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 0.714 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.639 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 45.177 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 159.97 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[97]
  PIN iot_out[96] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.61 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.775 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 99.9801 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 350.508 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[96]
  PIN iot_out[95] 
    ANTENNAPARTIALMETALAREA 11.307 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.5745 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.026 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.231 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 29.0929 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 104.327 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[95]
  PIN iot_out[94] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 10.948 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.458 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 84.9188 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 298.274 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[94]
  PIN iot_out[93] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.701 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.5935 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 21.1522 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 75.3201 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[93]
  PIN iot_out[92] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 7.908 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.678 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 59.6167 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 209.124 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[92]
  PIN iot_out[91] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.262 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.917 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 56.2115 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 197.417 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[91]
  PIN iot_out[90] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.004 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.014 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 57.763 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 202.847 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[90]
  PIN iot_out[89] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.801 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4435 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 14.8644 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 53.4035 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[89]
  PIN iot_out[88] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 4.692 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.562 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 34.1314 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 120.747 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[88]
  PIN iot_out[87] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.025 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.0875 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 60.1705 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 206.186 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[87]
  PIN iot_out[86] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.946 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.951 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 17.5447 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 62.1043 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[86]
  PIN iot_out[85] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 7.967 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.8845 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 62.9716 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 221.078 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[85]
  PIN iot_out[84] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.66 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.95 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 14.2696 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 51.1213 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[84]
  PIN iot_out[83] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.253 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8855 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 51.5596 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 173.319 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[83]
  PIN iot_out[82] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.046 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.301 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 59.3608 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 208.941 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[82]
  PIN iot_out[81] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.513 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9355 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 18.7344 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 67.1597 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[81]
  PIN iot_out[80] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.796 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.926 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 22.7441 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 80.7823 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[80]
  PIN iot_out[79] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.083 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2905 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 59.3198 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 199.999 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[79]
  PIN iot_out[78] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.38 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.33 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 57.9521 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 196.172 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[78]
  PIN iot_out[77] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.085 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2975 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 58.3523 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 197.693 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[77]
  PIN iot_out[76] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.22 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.77 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 13.7037 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 48.9009 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[76]
  PIN iot_out[75] 
    ANTENNAPARTIALMETALAREA 8.691 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.4185 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.354 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.379 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 27.9348 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 100.063 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[75]
  PIN iot_out[74] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.242 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.987 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 111.022 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 390.168 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[74]
  PIN iot_out[73] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 6.865 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.0275 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 85.559 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 300.744 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[73]
  PIN iot_out[72] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.606 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.261 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 19.3406 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 69.2816 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[72]
  PIN iot_out[71] 
    ANTENNAPARTIALMETALAREA 18.929 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 66.2515 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 7.384 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.124 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 69.1405 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 243.836 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[71]
  PIN iot_out[70] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 19.595 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 68.7225 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 152.384 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 527.809 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA23 ;
  END iot_out[70]
  PIN iot_out[69] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 18.849 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 66.1115 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.07 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.885 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 8.8191 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 32.4563 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[69]
  PIN iot_out[68] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 14.545 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 51.0475 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 110.226 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 382.537 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA23 ;
  END iot_out[68]
  PIN iot_out[67] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 12.867 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 45.1745 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 87.4804 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 305.878 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA23 ;
  END iot_out[67]
  PIN iot_out[66] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 12.24 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 42.84 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 83.7115 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 291.863 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[66]
  PIN iot_out[65] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 10.465 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.6275 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 69.2973 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 242.093 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[65]
  PIN iot_out[64] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 10.562 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 37.107 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 69.9296 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 245.219 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[64]
  PIN iot_out[63] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 8.625 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.1875 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 64.9208 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 221.332 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[63]
  PIN iot_out[62] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 8.854 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.129 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 58.7953 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 206.249 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[62]
  PIN iot_out[61] 
    ANTENNAPARTIALMETALAREA 9.613 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.6455 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 65.147 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 227.247 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.162 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.207 LAYER METAL3 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 72.722 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 254.672 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[61]
  PIN iot_out[60] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 9.216 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.396 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 61.1551 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 214.508 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[60]
  PIN iot_out[59] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 10.414 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.449 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 69.8889 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 243.963 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[59]
  PIN iot_out[58] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 6.445 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6975 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.978 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.563 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 17.8804 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 64.1708 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[58]
  PIN iot_out[57] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 9.302 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.697 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 61.7158 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 216.471 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[57]
  PIN iot_out[56] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 8.024 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.084 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.978 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.563 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 12.1069 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 43.7523 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[56]
  PIN iot_out[55] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 8.784 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.744 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 60.7285 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 211.536 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[55]
  PIN iot_out[54] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 7.094 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.969 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.886 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.241 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 17.3872 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 62.2334 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[54]
  PIN iot_out[53] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 8.122 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.427 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 54.9475 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 191.669 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[53]
  PIN iot_out[52] 
    ANTENNAPARTIALMETALAREA 7.519 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.3165 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.702 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.597 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 2.764 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.814 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 56.0183 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 199.267 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.94133 LAYER VIA45 ;
  END iot_out[52]
  PIN iot_out[51] 
    ANTENNAPARTIALMETALAREA 4.99 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.465 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.449 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.7115 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 11.752 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.272 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 87.19 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 307.151 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[51]
  PIN iot_out[50] 
    ANTENNAPARTIALMETALAREA 4.664 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.324 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.266 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.071 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 10.964 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.514 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 84.81 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 299.337 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[50]
  PIN iot_out[49] 
    ANTENNAPARTIALMETALAREA 0.064 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.224 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.358 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 16.006 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 56.161 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 111.377 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 392.11 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[49]
  PIN iot_out[48] 
    ANTENNAPARTIALMETALAREA 0.066 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.15 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 15.238 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 53.473 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 118.884 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 418.597 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[48]
  PIN iot_out[47] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 9.032 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.752 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 59.9557 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 210.31 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[47]
  PIN iot_out[46] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 7.292 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.662 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 50.5642 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 176.983 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[46]
  PIN iot_out[45] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 8.28 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.12 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 55.9775 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 196.186 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[45]
  PIN iot_out[44] 
    ANTENNAPARTIALMETALAREA 7.206 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.361 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.692 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.702 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 23.6698 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 84.9348 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[44]
  PIN iot_out[43] 
    ANTENNAPARTIALMETALAREA 6.229 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.8015 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.318 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.253 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 68.3739 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 240.366 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[43]
  PIN iot_out[42] 
    ANTENNAPARTIALMETALAREA 0.083 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2905 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 6.866 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.171 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 98.0238 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 344.673 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[42]
  PIN iot_out[41] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 9.152 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.172 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 62.1679 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 217.726 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[41]
  PIN iot_out[40] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 7.291 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.6585 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 50.4899 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 176.74 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[40]
  PIN iot_out[39] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 8.79 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.905 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 58.3781 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 204.789 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[39]
  PIN iot_out[38] 
    ANTENNAPARTIALMETALAREA 6.439 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.5365 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.58 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.31 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 72.8892 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 257.403 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[38]
  PIN iot_out[37] 
    ANTENNAPARTIALMETALAREA 7.642 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.747 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 12.424 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.764 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 85.1186 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 300.206 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[37]
  PIN iot_out[36] 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 7.456 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.236 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 54.8093 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 191.047 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.235332 LAYER VIA23 ;
  END iot_out[36]
  PIN iot_out[35] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.616 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 68.851 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 239.9 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[35]
  PIN iot_out[34] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 5.852 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.482 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 98.1157 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 343.07 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[34]
  PIN iot_out[33] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 6.581 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0335 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 105.205 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 368.035 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[33]
  PIN iot_out[32] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.318 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 93.2298 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 318.924 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[32]
  PIN iot_out[31] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.421 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.6135 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 58.8517 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 207.57 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[31]
  PIN iot_out[30] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.162 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.567 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 74.6659 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 261.432 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[30]
  PIN iot_out[29] 
    ANTENNAPARTIALMETALAREA 9.651 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.7785 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 9.6 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.74 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3328 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 55.4772 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 195.898 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.579138 LAYER VIA45 ;
  END iot_out[29]
  PIN iot_out[28] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.28 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.98 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 63.2396 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 221.917 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[28]
  PIN iot_out[27] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 3.919 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.8565 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 27.3915 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 97.4596 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[27]
  PIN iot_out[26] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.052 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.322 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 55.0143 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 193.928 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[26]
  PIN iot_out[25] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 7.953 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.9755 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 54.369 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 191.669 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[25]
  PIN iot_out[24] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 5.864 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.524 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 93.3934 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 327.022 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[24]
  PIN iot_out[23] 
    ANTENNAPARTIALMETALAREA 6.225 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7875 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 6.946 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 24.451 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 53.9045 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 190.756 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END iot_out[23]
  PIN iot_out[22] 
    ANTENNADIFFAREA 0.4012 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 6.624 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.464 LAYER METAL3 ;
  END iot_out[22]
  PIN iot_out[21] 
    ANTENNAPARTIALMETALAREA 7.349 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.7215 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.491 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 8.614 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 30.289 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 74.3035 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 262.819 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.94133 LAYER VIA56 ;
  END iot_out[21]
  PIN iot_out[20] 
    ANTENNAPARTIALMETALAREA 0.222 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 17.814 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 62.489 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 123.802 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 436.51 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.94133 LAYER VIA56 ;
  END iot_out[20]
  PIN iot_out[19] 
    ANTENNAPARTIALMETALAREA 0.249 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.491 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 17.262 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 60.557 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 120.228 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 419.512 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.94133 LAYER VIA56 ;
  END iot_out[19]
  PIN iot_out[18] 
    ANTENNAPARTIALMETALAREA 4.794 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.779 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.304 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 12.734 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 44.709 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 92.1829 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 326.055 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.94133 LAYER VIA56 ;
  END iot_out[18]
  PIN iot_out[17] 
    ANTENNAPARTIALMETALAREA 3.597 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.5895 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.3604 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 12.846 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 45.101 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 96.1216 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 335.138 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.94133 LAYER VIA56 ;
  END iot_out[17]
  PIN iot_out[16] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 13.274 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.459 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 92.7979 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 325.258 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[16]
  PIN iot_out[15] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.225 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 53.4632 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 179.994 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[15]
  PIN iot_out[14] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 5.936 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.776 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 57.6776 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 201.777 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[14]
  PIN iot_out[13] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 6.035 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.1225 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 56.6985 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 198.59 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[13]
  PIN iot_out[12] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.246 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 51.4619 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 172.722 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[12]
  PIN iot_out[11] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 5.865 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.5275 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 56.9645 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 199.161 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[11]
  PIN iot_out[10] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 6.148 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.518 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 54.559 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 190.735 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[10]
  PIN iot_out[9] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 7.545 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.6875 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 59.6789 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 211.076 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[9]
  PIN iot_out[8] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 7.12 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.06 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 54.836 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 193.516 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[8]
  PIN iot_out[7] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.281 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9835 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 66.4358 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 225.385 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA34 ;
  END iot_out[7]
  PIN iot_out[6] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.462 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.757 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 19.469 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 69.1995 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[6]
  PIN iot_out[5] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.085 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2975 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 38.7793 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 135.939 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[5]
  PIN iot_out[4] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 5.832 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.412 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 81.4977 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 283.967 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[4]
  PIN iot_out[3] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.503 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7605 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 40.9593 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 143.689 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[3]
  PIN iot_out[2] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.694 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.429 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 45.7533 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 160.014 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[2]
  PIN iot_out[1] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 7.775 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.2125 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 95.4443 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 334.08 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[1]
  PIN iot_out[0] 
    ANTENNADIFFAREA 0.3604 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 9.908 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.678 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 123.521 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 432.349 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA34 ;
  END iot_out[0]
  PIN clk 
    ANTENNAPARTIALMETALAREA 0.09 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.15 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 18.754 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 65.779 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0754 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 503.552 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1767.06 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.43634 LAYER VIA45 ;
  END clk
  PIN rst 
    ANTENNAPARTIALMETALAREA 6.33 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.155 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3952 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 26.3529 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 89.5997 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.0913462 LAYER VIA23 ;
  END rst
  PIN in_en 
    ANTENNAPARTIALMETALAREA 5.589 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.5615 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 22.956 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.486 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 21.683 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 76.0305 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.481 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 68.3854 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 241.018 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.705997 LAYER VIA45 ;
  END in_en
  PIN busy 
    ANTENNAPARTIALMETALAREA 0.062 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.217 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.886 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.241 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.3646 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 13.854 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 48.629 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0845 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 184.341 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 647.711 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.28166 LAYER VIA45 ;
  END busy
  PIN valid 
    ANTENNADIFFAREA 0.3604 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 7.008 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 107.801 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 375.994 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.544495 LAYER VIA23 ;
  END valid
END IOTDF

END LIBRARY
