/opt/Design_kit/CBDK_IC_Contest_v2.5/SOCE/lef/antenna_8.lef