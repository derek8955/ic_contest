/opt/Design_kit/CBDK_IC_Contest_v2.5/SOCE/lef/tsmc13fsg_8lm_cic.lef