

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO ISE 
  PIN image_in_index[4] 
    ANTENNAPARTIALMETALAREA 6.568 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.988 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.002 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.647 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 44.726 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 156.681 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 2.436 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.666 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 112.552 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 408.839 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 4.20746 LAYER VIA67 ;
  END image_in_index[4]
  PIN image_in_index[3] 
    ANTENNAPARTIALMETALAREA 6.732 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.562 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 8.88 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.22 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 41.468 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 145.278 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 2.436 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.666 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 152.552 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 548.839 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 4.20746 LAYER VIA67 ;
  END image_in_index[3]
  PIN image_in_index[2] 
    ANTENNAPARTIALMETALAREA 7.47 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.145 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 16.332 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.302 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 42.88 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 150.22 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 2.436 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.666 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 188.823 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 675.786 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 4.20746 LAYER VIA67 ;
  END image_in_index[2]
  PIN image_in_index[1] 
    ANTENNAPARTIALMETALAREA 6.322 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.127 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 23.692 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 83.062 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 42.522 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 148.967 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 2.436 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.666 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 224.627 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 801.1 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 4.20746 LAYER VIA67 ;
  END image_in_index[1]
  PIN image_in_index[0] 
    ANTENNAPARTIALMETALAREA 7.224 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.284 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 33.628 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 117.838 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 41.436 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 145.166 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 2.436 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.666 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 150.921 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 543.128 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 4.20746 LAYER VIA67 ;
  END image_in_index[0]
  PIN pixel_in[23] 
    ANTENNAPARTIALMETALAREA 6.978 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.423 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 23.784 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 83.384 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 16.548 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 58.058 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3588 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 76.9706 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 271.767 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.09615 LAYER VIA45 ;
  END pixel_in[23]
  PIN pixel_in[22] 
    ANTENNAPARTIALMETALAREA 6.65 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.275 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 29.58 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 103.67 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 16.334 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 57.309 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3588 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 64.6208 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 227.809 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.831382 LAYER VIA45 ;
  END pixel_in[22]
  PIN pixel_in[21] 
    ANTENNAPARTIALMETALAREA 7.552 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.432 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 35.294 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 123.669 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 15.146 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 53.151 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7449 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 39.6131 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 139.218 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.750444 LAYER VIA45 ;
  END pixel_in[21]
  PIN pixel_in[20] 
    ANTENNAPARTIALMETALAREA 36.496 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 127.736 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 49.462 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 173.257 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3679 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 143.889 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 505.429 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.800106 LAYER VIA45 ;
  END pixel_in[20]
  PIN pixel_in[19] 
    ANTENNAPARTIALMETALAREA 34.402 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 120.407 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 38.638 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 135.373 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5525 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 80.4349 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 281.73 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.573864 LAYER VIA45 ;
  END pixel_in[19]
  PIN pixel_in[18] 
    ANTENNAPARTIALMETALAREA 14.774 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.709 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 15.524 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 54.474 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 21.218 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 74.403 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.663 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 65.1923 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 229.083 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.1506 LAYER VIA56 ;
  END pixel_in[18]
  PIN pixel_in[17] 
    ANTENNAPARTIALMETALAREA 13.383 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.8405 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 21.602 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 75.747 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 21.3 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 74.69 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5538 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 54.1784 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 190.471 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.701455 LAYER VIA56 ;
  END pixel_in[17]
  PIN pixel_in[16] 
    ANTENNAPARTIALMETALAREA 7.608 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.628 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.042 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.787 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 26.37 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 92.435 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.572 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 73.403 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 258.322 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.596889 LAYER VIA56 ;
  END pixel_in[16]
  PIN pixel_in[15] 
    ANTENNAPARTIALMETALAREA 10.256 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.896 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.304 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 23.392 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 82.152 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.351 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 95.1496 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 336.2 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.199 LAYER VIA56 ;
  END pixel_in[15]
  PIN pixel_in[14] 
    ANTENNAPARTIALMETALAREA 7.332 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.662 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.714 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.639 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 27.198 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 95.333 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.351 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 102.622 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 361.953 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.199 LAYER VIA56 ;
  END pixel_in[14]
  PIN pixel_in[13] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.98 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.796 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.926 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 36.49 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 127.855 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6188 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 77.078 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 269.923 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.847447 LAYER VIA56 ;
  END pixel_in[13]
  PIN pixel_in[12] 
    ANTENNAPARTIALMETALAREA 27.406 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 95.921 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 14.654 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 51.429 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3679 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 74.0773 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 259.089 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.561634 LAYER VIA45 ;
  END pixel_in[12]
  PIN pixel_in[11] 
    ANTENNAPARTIALMETALAREA 36.22 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 126.77 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 25.72 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 90.3 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5525 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 61.0925 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 215.058 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.06737 LAYER VIA45 ;
  END pixel_in[11]
  PIN pixel_in[10] 
    ANTENNAPARTIALMETALAREA 36.17 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 126.595 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 19.492 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 68.362 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.142 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.137 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 17.609 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 61.7715 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.663 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 50.2453 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 177.179 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.839668 LAYER VIA56 ;
  END pixel_in[10]
  PIN pixel_in[9] 
    ANTENNAPARTIALMETALAREA 7.306 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.571 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 28.834 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.059 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 35.328 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 123.788 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.702 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.597 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4667 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 17.3635 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 62.4794 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.976419 LAYER VIA56 ;
  END pixel_in[9]
  PIN pixel_in[8] 
    ANTENNAPARTIALMETALAREA 7.47 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.145 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 18.458 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.743 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 30.1 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 105.49 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 2.726 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.681 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3874 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 24.1177 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 85.4103 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.514888 LAYER VIA56 ;
  END pixel_in[8]
  PIN pixel_in[7] 
    ANTENNAPARTIALMETALAREA 8.29 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.015 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.806 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.461 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 27.896 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 97.776 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 5.486 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.341 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 43.8763 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 153.008 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.03775 LAYER VIA56 ;
  END pixel_in[7]
  PIN pixel_in[6] 
    ANTENNAPARTIALMETALAREA 5.912 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.692 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.426 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.631 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 43.034 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 150.759 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8554 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 57.966 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 202.966 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.772972 LAYER VIA45 ;
  END pixel_in[6]
  PIN pixel_in[5] 
    ANTENNAPARTIALMETALAREA 5.912 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.692 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.426 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.631 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 12.604 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 44.254 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.334 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.309 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 18.036 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 63.266 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2522 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 129.652 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 454.879 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 0.937946 LAYER VIA67 ;
  END pixel_in[5]
  PIN pixel_in[4] 
    ANTENNAPARTIALMETALAREA 5.83 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.405 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.334 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.309 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 25.61 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 89.775 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 7.694 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 27.069 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5902 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 67.2823 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 235.834 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.26376 LAYER VIA56 ;
  END pixel_in[4]
  PIN pixel_in[3] 
    ANTENNAPARTIALMETALAREA 7.224 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.284 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 12.192 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.812 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 40.676 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 142.506 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5694 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 91.5701 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 321.55 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.794169 LAYER VIA45 ;
  END pixel_in[3]
  PIN pixel_in[2] 
    ANTENNAPARTIALMETALAREA 6.322 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.127 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 15.596 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.726 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 33.04 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 115.78 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 8.797 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 30.9295 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2522 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 79.3971 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 279.82 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.01705 LAYER VIA56 ;
  END pixel_in[2]
  PIN pixel_in[1] 
    ANTENNAPARTIALMETALAREA 6.076 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.266 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 22.598 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 79.233 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 33.39 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 117.005 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 10.249 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 36.0115 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6162 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 41.8966 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 146.684 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.847939 LAYER VIA56 ;
  END pixel_in[1]
  PIN pixel_in[0] 
    ANTENNAPARTIALMETALAREA 9.079 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.7765 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 41.652 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 145.922 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 19.838 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 69.573 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7254 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 46.0014 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 161.903 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.52675 LAYER VIA56 ;
  END pixel_in[0]
  PIN color_index[1] 
    ANTENNAPARTIALMETALAREA 7.976 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.916 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.026 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.231 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 3.2232 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 48.777 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 170.859 LAYER METAL5 ;
  END color_index[1]
  PIN color_index[0] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.98 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.174 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.249 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 3.2232 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 56.894 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 199.269 LAYER METAL5 ;
  END color_index[0]
  PIN image_out_index[4] 
    ANTENNAPARTIALMETALAREA 8.712 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.492 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 19.696 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 69.076 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 3.2232 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 46.089 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 161.452 LAYER METAL5 ;
  END image_out_index[4]
  PIN image_out_index[3] 
    ANTENNAPARTIALMETALAREA 7.792 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.272 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 28.132 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 98.602 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 24.622 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 86.317 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNADIFFAREA 3.2232 LAYER METAL6 ; 
    ANTENNAPARTIALMETALAREA 3.666 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 12.971 LAYER METAL6 ;
  END image_out_index[3]
  PIN image_out_index[2] 
    ANTENNAPARTIALMETALAREA 8.16 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.56 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 39.796 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 139.426 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 3.2232 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 50.086 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 175.441 LAYER METAL5 ;
  END image_out_index[2]
  PIN image_out_index[1] 
    ANTENNAPARTIALMETALAREA 9.448 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.068 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 44.972 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 157.542 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 3.2232 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 47.99 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 168.105 LAYER METAL5 ;
  END image_out_index[1]
  PIN image_out_index[0] 
    ANTENNAPARTIALMETALAREA 21.776 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.216 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 50.588 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 177.198 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 3.2232 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 3.83 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.545 LAYER METAL5 ;
  END image_out_index[0]
  PIN clk 
    ANTENNAPARTIALMETALAREA 0.254 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.889 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 28.016 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 98.196 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 49.176 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 172.256 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.3 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.33 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0754 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 33.7115 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 126.329 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.91512 LAYER VIA56 ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 14.88 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 52.08 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 28.266 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 99.071 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 332.848 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1169 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.02849 LAYER VIA45 ;
  END reset
  PIN busy 
    ANTENNAPARTIALMETALAREA 61.572 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 215.502 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 3.2232 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 22.444 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 78.694 LAYER METAL4 ;
  END busy
  PIN out_valid 
    ANTENNAPARTIALMETALAREA 8.886 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.101 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 13.382 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 46.977 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 3.2232 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 52.037 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 182.269 LAYER METAL5 ;
  END out_valid
END ISE

END LIBRARY
